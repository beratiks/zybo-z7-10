

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Oz3bq1Y3q/0V9ixcuZbHLMVuCmNW1UJyldjpAI7CeoQPTqDZudIgrgjWR9NF0qCtBLJSCMXzP1Sr
eN9C8zv4sA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KWRaLoIwCsXaL39b9IKN01JCLrps/lNaWQ7nl3x6ncUNUlhw/8FEb4bwWUu4OR8OSSzcmb49sqFg
iD+mFiPB/MBPMZqORtlzHg4I8jIpTQLqgrFoaXNGaz8egy2VgBuHLge8oxc9DgFyx+QRrX++gBQo
zKjdvnUyXg42AfFbvEs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
1IEFoMViZkns8aGwNXB0xHaJtjPilfH4hlkwv5gIB4hPzjNJyT9JVdow2VvbjvAduNrsA9FAv80v
G8Q8RP9825geM8Zi2YxrJTgHodm6Z2zBVNgCztCtQGXpRbaCmFBL/zrjjOjFKLXIHWDYQLUx1kcX
e3rhReJ+F7v63rjet5zZa5OZ8ogQHdR2nzNNpbvejOJ8jsY6ZjfboXTwo2/jzRcV0K2L6vosAuUW
A2NfpV3bz0zFVsCIAd13ZJ9T3sj+nO3OsbDV5SOHm2Ren2bFJcjgVVtLMgDtdYUUdz5BrMreid4D
zCW84ekERCzzZD2EtVZSjHAg1qKpo7OZ4Ou93w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Al4qgSgowgaB7wG2rIY9SCMsPkMatdGRWZ+7S6JiJvwZYY9+OGBfE9b6SOjMAb9B/rD381e63NWR
SDfChuWksMWI6gFasoLRMRhek2eHqqGaTg0bmxxbwNqX/7UK9581kco9v68YfdVceyETwNKCMSKX
e4hryAFWb9CLPvGXeZ7mLgaAG1VOjoBtolhlMPm1hwiVrDmdeiVAxP1xPuMDZCp61+Lb6j1ZsiaN
WvVdmJEZS1Mk4UuwBfWw/Ch7qyULfDfcISPKjFv4sm7FPXpVgb9ajOHjO5F3i67qUFYcVt65UgC3
71X3EN/lSdIfI7pRoSCLuH/clQ7prL4fDB3xLg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AluE9BIse3ig/Scm50r30ADy/v4PwTkEbRoIJ3d1ekSZO38Oc8kFGVvK7XJWDEffYBXKxMz1CccA
7BKnsot4wFC8u7cmjnltSZVWQP47VV5fjw+gMZ0iHULvWuRBEeAKtgBM7ykDGAIUJ7V6klpAAffn
a2wgqu9XC1kYHN7+vcQp3OSFnlTnFFYHEUWVgSo13IOa6dfcL+jxSPVjcfxBsjz0dbC/gkMbDLZl
R2G8+cnZgvk96wa9jv1r9MjNzZ1q+IwL8ASXqrsI0yPd/YZEmCvq1Ny/SeoxQQKaRejyNoO/NsB8
oIfGKPVHyn/NhOlXciQRtDFoVZuiIucs2wTLow==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AR2vy4QzCevoZ+e0bg5vysvbM4wHmPo+GktognNJYBUj5lqIeHWmOxyP9yhgLiqeFoLBabBOo+Iv
WtceE+75LMJBYUiYjvS9oSX36qF3UWrnT/FxFG5xEtyDeNyFC6sZ78WNMgwqptiPGhNYwy9Doh+h
+ymTucPIk4JobvLKL+Q=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ab0HqEC7etg4Wk8pCsdzqJKhZFczgrIsDzDfy69niLkPxpIb+twU2iUyNOofId4FbKPpoDsA1Rbo
WChSzWh6JCQ6/gD0VI/tqImGVY1stdbfXfGykVKr8JjVy3BIPwuSeZQPhff5YRY3pxiTzpS6Oc8y
l0G3gFLO94CpFbaNjGijADVhLi95R7pu90WzAmQN7CRdbH4SmtpoXggdHOkugLGwsc+xah5O3Mqt
UT3GV1ppBSc2OMqUOzoaKe5iJP5QQgn/fHrLeZGxQsB2ha7xenSodqlX6ZCx5ZXhpaxi/4oNN3cr
DVTSNKSg45LNcntctf4IK99VIcUqbViGmn+lsA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 710400)
`protect data_block
4PGJ9Q+6GUKbARZinx1T628d/8HWjH9H4hcXkMw+sxcA2zrl2a77MvscnWC2ElAOo/LQq9Ciep4W
vWirnm4YIvTlrkk362loYx9i+gkTbh7PUD0abohIZe49mnK3pNdVAbFXRoaW+8XUoTIx90uvli+K
bafPN+yqvaPdpVKwuM0XVyipHenUAvyk9qbIGN+PRWmVsBthOMslt2etY1HxtISjg/NUhP3qJLhC
GeHQJZyrmsREEEce79bd7W3WBlIk4ARO5EsVr2DzP/bnu6vtOxiYOdgGHj8LG/Vv6Tm3m7a8u55v
CNgNW6rycIalhs4rYZ7zkQ68PoIoi5Q2GuuGw0sHLRxzLpBWTYMruJP98TqQYQRl9yO5pGPrKeDL
4YEK17mjAAfjllsf3u5z0jLShZaQbibwobu5GTNXcibUbfRxxrfnSLMm9tHIzqqwr0tWHNZdntsw
iH2/drTRlTJ8Cx6wPgPNTL3OFSt84rDFyTiVdXBYEHU30MXt1PLsRp2FyXu0TIq/eEm6muwYV59j
w5uh8Yanneq3XS3EOp6dDOMy33bbX12ITCz8sWoSVXCwJQZap97hxrRYwHYRCBcqSB9vaQEpOJE3
Xcb7xf44k3t+LbT6cnDjJYX7vOdqdXBb245TnKBC8bCU97QQ1OUc1QV1yx8nms1K9lFRkEs9+QLA
XJW5pPcDlNvCpQxklPCXprSv8moSV91c2S9SmzVUJIrdSB9L4cmto7OhGtY0E9GkWt9ELatLWY1Y
LvA+o5THGPHl5Jkm4sLRJsPA9l+ghdbNIzHfN/sKYpVuE5HhOO1K4pp2LAMeCaaFRAGsWlwiwRnI
tvjnVLJlx1ygZApQvymho9+Y2FoNDi9MSPVmQa+mC5uiHx3Qx7zV5qHXcUiNzMuUtf7x3km5LeSk
71+JjpwHDJHBqGjih20fph8OdPvHjztQKLtEE5t1EpOgQXRBW899l//CM1KbHlWd3NGlaMOVeCQm
JeWnZlIY2XrKv/lhx8ek7cVFfQkoZnpLgVCPtJfYKmsMoF855Uo4Qer0hbgVfCoPcadwbU9uYNcW
T7rztDc81q+06hTuXPtIK/vHxEaJWiYdyVjmuzOAWu8jhOA07XV3QDtlYaHD164Wv+fQuDJdk21U
5f4woCGhCao7mTeW+ME8ccb9k0R56XQbwhy34b19LJ9WJfkGoy7xTTlV/Wd2R/dpqEoASl8gi+KF
d4YP4m9laZ8iwb4wuH25TnWY5r0ig7KdUk3dGGeM8CCmF5tcznFz1WCM8RZWVdEK3/6NErG3coFr
B8N9986IvHJlL22TmbJHMgW0njrHGpz7RKepWkSQkoXiY3PzLCuruVih4WqbnaXixKz6mV0urC2e
tz04fo+X6BopPgv+i/S1av4yza0p50kjjoHqo2e11Lga+bfEnvPgQL2exfTtfbspq+7CLETiw9n8
3pFU2lW4jwnyIAmwG/eI7u5UOzI1shJ8RG4ORUrKl1fYPijEtktLP/36V/8qbWcAN8VvxYtwKADC
MrLHro30liVHH7Rhxy82q30rQf854lXe5PLUljCT2n3bs2Ea+arFm2y8a3suVwSKmeTklm8oSt1B
Ezd5F96sX6yb/m4/4+h0FPDssgpgkE4u52G0ssOHmXNolPZ0QKWJSd9wC1Ta1PNuLpDtdSdD1O7L
kgacpjMwVhL+EFG07IXmON+rqs8pO+VpsVa2cRGE3+mnbzbVxNe0Jr07AmcJpK2+w4+6weKfdyNR
tuERdkqq5NELpA6jDxLqDZXhvupA/WPVmftBt3Rbb5lLVbY9ddFhvIbR4ivCSE5qknqzXVZv6IEZ
KUVMUt4bqn+aprZTnQ5h6TmCmHWklqPtnrDB0axNhuH2oHOqnkvxtDjKWUDy4V+Stieb3bz0MlZk
f0MlTNPgbuIanVSN75+MUnwILGixHkP0rX0owpyTT1SUrznLAXSz8/JP6WjN3jztOMCYOqFbgImt
OF/d/BIK+dvl/Q5x3CmXwLy+GIgThuT1xuI/rldgWLyK8ZJIy2eegulwKLHsfex462JaDvwan8Wn
PbkZaabDJYpnnWvRS+EBpkbc31fdtEXvsLiTcsiTsVFpjpXCvOwguGjTqrRXp99FzW0pBMdIfr5W
liqiDTSj6S1gydlQE2nlQk39wLpG5Cy20dbLwXMQjHl3M5c6V1Lv6hcIXKlZiQ+GwGL/EpmoC9ws
cCgtGFl4NsCEDJcVBeiu7Ene1tUXn6yEMz0g/gu/kcSBFGKNHM+9cDRmWE5wCpVTuMVBRxeXbrFw
VxjFLoxVm/kBPdmXi20C3Wcn+OnRTxft9bp6mSocbk4fh56bNekc63vKUj7hVVNGcwz1YkX2QAqg
MwuVrIY40re4gFAf+OTHkECDP0eQ1DCD8TIr8+YgKUpu7itBIyhJaqFAVA9bcyOBMupRLDLEWj/4
k6yFyftuwb6Nb9aYQgso14Bx9Kg8bHnuY5q1bDAGXhIdS8YMXUEFePi+omT7Ig9E6FzMdg2dUJCY
vbCBIpK7Uf2cx4GGkb9NLRQm/EiyDvk4KXD4nV1iVrqrXIdLsJG5fdt1mFvlt+EP6cqtndj1IGrO
piLu2xHvIpm8knGIjKC7upS6TxNr5BtVmEx2+gWZ1vt3wpG6wADqoQRf3/VuiD5AfkhaSi5i4+Fh
zKYfCxUqJDUcTVDCWxdkjjxMdPinncruUQI5sI5gAC+vXKxw3n2oIfSANtpdm3okbKUHIifiaSLx
+ZdMxOsz/oHRlOFslePGSMWyV5bD0yS7FRBwJTEgZpX1bqWXKf5k4lokMLBY9q3YHFa3YZRaHVA/
p2g/y3eawsdpa9lCE+qZNlsuKI35lxljy1W6zt1AI66RKn/F2zNKDBwLhAbMhuSy2puh/JnRIcOi
BW5zbPRF0HxN+9UCjhYDIg1NXKXKGiJI+nwTdrZACSGfYJLF/SB9eCnyXpRcjW2pVI/E4RcKR1SI
InqlbJqYssIHhdHC6OAfpJxouMGUXk+0yj4UTaVJIjBZBuznGf2n7qxwctESxgM7LP5oxN/N74vz
z6lBI8xXsemEKE/2VH0Q6YpOgDaEHyFHPtmqED8ow+GCh53p6D24wz8dxytXk0hT8p1Z4YPJzT/m
QuDfZTYIpojgEVm3OD80Y53UH2JZP8edIz8ypY2x36pJgJOSt1BMFqYbKFrYmRFb5H91A5uvpDwJ
8yPCkBH+578ot40UDnY+K9CTXh0PRlEfI8SS730v4Qw4FHhFuFjuSL7pZuOhtiSO85BUjTrtFrxB
XsqSL2qG0JZJXXlQ8QQXtj6wYzure2FEakXwFqYBeKUZfQMrkyMUkZKusvl8+X9c3MvaBq+RrAOA
FYj9hbCYPbhjVrVr8Aqj/O+ZaUv+gk1ZzTJ096NquIUIWAHkr0r4k8aQJKr6QS2fu3zqp6Qonp/m
RPNnfDp3HpUyryKJL4lhjRvuRACHqnI1+xkazmDa2oMcjw8i4znEwQXo4sv4YuWxW72zVH9lpOiX
Y+PAYFWpLx+BKG7jXpsYpdk/JPj7fd2/HZ0GnqxvVB7NHpOVGC2TgyG6x7x+z+61S5grdzVZ1/rB
4MUdSVbK4udIq4ZWoSxiHhJKr7zdwbvTk2avpbwfaG+kGYoDq6D8plkeb/9L4dLKeYAb852ySvxj
i89hHMOG9a+3cOERYS0NPx8BAlmB44wcHmAX+IQ5YOU19cENy1Hy1+NsLGqldHSS3dOGXoEYM52S
FIC7/bDDP8wnMUWuDUzK+IlvRnW0r183xFguboUpMXxTSs+pdurkbstZbY/BKc/a60nQHqZOWVf8
ib3GEc7Uw/Pym/WIl8Clm93r5/5qMVIoCQ/HBxEL91J6cXCdJrStHzWyVasn1UchxR0OlpdKttKE
//4aHdnQ4H1eee5tkEvYpurgVO3BqxQHuzMZiSxAGRHRKYbXfqH6NsC17odo9uyCiGvkE61ITFrV
q6wjFFGZPLaztuNBgGY14n+6U4KF+pucxFHa6IqxGKYOIYbk1aDE1rEX2UFcNY1abB1VWfPLtrwG
xMQdsCrIrUxYp8S6IOz576g//tNpogSr8m792ZzqxVksPqsAUG1xTgS2y8YBP0g5Wfb3itSX3sv6
DiHmEPPvsx9u80tHmSonH+SZ4iRO778PLZ6lBlNxZA86I3kk6jiPjhvxJB70/5Kd0pPKWk8E9l51
Q3fdjWQesi6FRQvvTkGZRXX+tvlW1LPFj56H4FseqeMlPIPCv4thmUxWGdy7fmWdXUU7dXF9NugK
9jCDyuAYM35dw1GlsT7fwJeLS3Sxo3LnfQrBSxh8TqRY8Zk1E9bBBhCCF4qKauGnrnJdDAmyhc1g
3yizBLuAOKPfusxbXslALOPCPrrObtwPA4UZCQspPi98FfAL8cPXbbykl7cftdEAYdkMq2oOdorF
9xN3jDahr9SnfzbVqzAy3w1aNJyZ1x3+vyVUcXE2vMIGKh4Y/G/RHp4kfkVvO2MCloKlx+8YAjWl
Aj2OTWut1Kml3WFehzvPXktflir4vmU7RmQuMTURCztts7rJbSqx9qC0U5qkGuXlPJvBunD3b5C6
0O7nBvWe1vW8PlAJW2A1GrzIi0vuRIjZShptHygBUE5A/jDJTV53oP1pG4xW9/+akVYwFSoq5lDt
W083Zgl3xhFkG5XY0+p3QLAyw3Qz2lP+pLCVWouyuKUqEsoERyN+zGDys0MV+4uuHieVr55STasO
OKcg1oRYHVluj8N+kZMaUfDDY5W1RgjBSwTkEl22oNv3gH89ogH+vgLxCgxxnDFXq6oN1Pg+0CdO
q9gjrCopwsNh3860oLUCX/rcgrnys7YrAAS0r1NqBRI8znCQnmyXXMojef4PdB9MjHvAXmN5rY7E
R/3gIkj20T7E+TtfeDEVbod2OKjXbIHnD9cKi19NcbTUrDP5beCNV96K09kstEKYTRYeelYO9qsA
mPnvfzyC9oFSOYAd2aijLzGYgQ53/WuMwuMVDEcWdmkCJ9ZIsH7oStBiUD0bSSs6gYU5JOKnbkKa
JISYXEHHbZ6mfqvA09hyQcyFbXR52qUL82y6fYhHyZ2sWa88qZoZ/yPZIDPmiab3Vw2htQdc2p/P
ZVzLiXhHvu+PmZbDA9uPNCJ7L2sIU9B3n/f3Qco8yFeiL07H1O/nzmoIvKChPXALXI1sclnwu7cC
yzqOrzSc1d2w8bj5kbclhK7yHww6K3GLGQBCwK41eRWNHoB7JyJDy8ymVwbrYlkFe/zgGEJGSg5T
RGjUj7SNrNtPxz4hlBe6/fQI4967nMLNvsPrIP/DdtHDgWY23czfNgkK8eM7iYMcE7Jxyug39X2b
7BIQXSCpaMn9ntw618fRqbUj9PQOsyMHzTQaZ9FtvQCTI3i8BJNyCBinKUG/CMlWU8pqiVKddKd3
9QuNLjppijiRo1bW/9UpknjLCLtK4YFf399Sb/zTZAegC4ZkRrTwLkXafD6SKIjABi4gT/IHuj1u
5kenwQca4X3KR6n62qpxyMcnNcce6Imhp7wAE4+tufyILT1tVtt1JbxFvxeDqzr2pQdPy5oWW+sS
t+Ust2gxizkitGTq2XEcu4H/644jflHPI9F0aQGT8N0zsqL5d8PIaQtJOs7t6YZvdsm8xsN0J5JP
dLPOI0ooDSnA+txOgLdlVdkrMMmloadYTXUqjkRbyQNenSA2Nbo5bIQXDsrKX3Q3gj9QyU+7dzB4
sNr/M913oHDdDUye6pjiHnBQ+a/XLxB5JiSRj8qScEgbTu78wGw67NWKC/9DbtimvASKGNNh6f+U
aKA13fSlU/RcB9H/LFI0pNuL8kuoHAglyq1YyukTV9w3f8c/Z6qylHM/YrZhRBPl3P8OiDe76onZ
aXIlh6+X2jiRMWZsKVLak6Cb9RGjWgj93IsVsAVGoguAGWf/xQ2TZIJcbt2l5k4SMGdJ9OtSzYL4
nOhhvcVWHQW15hU7u2icRLs5WmtvNa0K7YKFBikc+qjB3mV20bhk2p8zTh0vGcmz86m7hkIEuMvV
h5wE+kgdX6vkFb4Es2iyO5gfA/qg8tbZE0p3ozTUGUskuOxXlBlPy3vUr7O94EXxgJU9v+2qg7rQ
Vl/J7+zpFianrNJJs88HEVEIInsOwD//u1w+T6UhCDM+x5zY9GvKczolFAuZpw8cZ4IKIbV0IsvV
r165uCVOku3fByOLOXb83N7jhlIO/cA1XAU1INqccss+Oe+87djWqud/0Y83MuROgtht0y9c56qi
Prj6+2DK/bzE683HdeiyK45fuUB6KwzIOsuaaLhgoUkyhwRQkKBHKFcJj/TMuLvG7lNfSQasYWE+
n1V0NQqqGDZtpD+tb546jug+FLc4687cYqI1Jy63Lk3bIWQuggIIwMTb8SRsVsKXxSJgykpTAmnV
zouQ1yZEujbhmETQIlXc1zSz4PL7NvbTN1RQ9Am/KQbmC/aXwIYfriWtyK+fJ3eAuKxzHChC5Ay7
KOzDaPe56vUDbOl8JMEgEGz8OuBrql27FWCquDH2YG6NfWQWYmrt/FzRLycsFC3Bui/Wp3t7pOTu
YT5ivu4058uq0elT5ZCuAgRi2KhuViy7hALp07Y5HsHj0IrcAHPDD/1uDNCjnlUcbat2AprM74R8
0DS7w9oITHlW56z9tGmSYIthCRW3OOZ3gyHPh/VIWp2SHFB1cG7LLeVMFEZrc044Q+6tHaB/bB1E
pJthttboqXqDi7cTn4l6KuTNC7b510VciRlZg6HLg6ntiFatJf/mzLy5l0/0TQxQUZESLIWXBPdq
7TRX62V74k+RkdODDMZcmlVSo6SsA5NGRhpOqLflGWwAH0UlL4pdFKFtwhFSUHeQWorWBZGF/qBw
iISIy8vxF2jdKXzwWx/nwexwGdl70V70XSC/KVgD7/CzLxKPTShLZv+guQRBS0ck7ZDTP4LEJ173
Ls7ECqkEK3w7mx76spODjRcnMt0WOl9LrFKg5Xq9M7VQdlIG5nAUD5t6yjg699yJB8juIganQyP7
zGcn+jW8b6mn3rcw1CeGqcZr5NW1TUM0FZZsoo20c+2XQxm64lQ5/VMp5TEjptYaRCyKOqMp/pi7
1hTNOnCubRxJvYbrAio1AFXjCWSpHRlBQ1CPjdvQcDid7KLReJO5rCU0G7ww53NjT+nNGaAJ7Zy6
Wt0QgEWw0P/YORlMFfwI9bl5dBQfS2QxrfLW8o4AA9+/879GKvRkXs45SAFUase84nCRM0IUNKl1
1m0FM9OE6LQfxbHrSNd02zzy4WFcd2zhUedps1T3eFLP3AliBogfiEgnWSJ1BLk02qWqEKzRsJPY
hXQBQgI3CYUenBxuidcqq5mkXujX/VH6GkIx/P/6vRHHSvbpNKgHJ63pQr68JvdFWJnu6caq+Vee
UpxFBeo+lcSPQ/O0sSyPazzZk4w7rRD3V5rY/fHPijb0DVVOziTAHZnMbLvCgH50e0X6soQAnND9
ICHT9rxMAqt+C5DijeYPJ3UQltP1Vud9u8UcxAMpnqBWPhweSE9zvwQ9UGaFIfSh1mMwxw/9TnPd
xBKF18W+t1Y8Rd9VafIscVwwZZZM/qACu+akm5mI5tUrjzc/Y142AO/yKQep7j9agXDiEAYS6+BJ
2xlblZsXOU2Fxs52/sM7/Q5tBGmSrPQwu/q/2/Ljq1xhCTSuvTwhEMO7mRJ6OAyRvLTBPnLe2VV/
Cy6HsilMQVf/WjFVjdY436QTfog3bT3jMQAwFFZQ4I71zc5Muqcu8oQ4HvRbVTDPJEJt4z2c8d4O
VGPF8IDTAn1FFd1A8Ga1fz0LxFkubFcG2+KPN369Y6/YTg52Gd1lPVavCQv9BSOs2PGEDAr+utAE
8i9w29WzXHkfv3vOpsvLJRT2nGmdFQUZTYjXC88GU0ekKuviJBIp/wy3I8umnl0DJU76NK1KRFCk
lYqZy0dAJfH9GmDucCDIJjTMZbx6fDcZooQmkabPcjt4jGiWAWaqeY/vwY+CdXE0TIwpfC6ncpcW
TD49QXfc9dkZd+pKDDUCANzW/HQ1ifEjjN7zuU5bi0OZCtrS2gvoqA2zdMYzexQ4/Ox3nhHkeBKi
4P27D3CeLc2O3MMcfzcaGOxwqFnSRpOmYj1Zl/1yEvknZQZvQM8EPFBM32P+cgXc78SKEHTLGDpc
O9udrXRQvOSQT/bSGombOTNB6xYeXl1BPNP1BHezg96B4F/y8MJwGtO8Ft6ugcJutoxHNH1WSXol
IxQUK02It0GaDbXbdGt//SzrcbTCPcwB7YibkX/SPzJ52a23TAvWlBIzu1pp67V71hWJ90n/LUdZ
8MK+/AQd/aM+T/6QP7/+aCIGjvPdV1+10cKc11DJz10fzzPYwKBvY+LFXBj9Hh8+/yA91KTcWEWB
WmM42BYfxISLnIDzJuG4AydEGfdI0Pm0JFajtZN4LCq7JhbzzH0wD00rK367O1lH4FbOa5KALaPp
5VuTVJmCCwOJ8whtil/xL86GRRpWAOHHu7ZeCplyZbHKlUHYwLU7iEAsLg7VXRNJ0HJFu46lClnz
7Tx+X5yGgQU+o0Fav+FsvM+aSS78IXG4nYOgTf2hCrRbSSuzC4++UdAlNjoHKDVM5KnE9gpeidpf
qv6u2tJBcoBTixcgO+hRmvNUHP8fzundJTe/hmOj2bbZvllDak6IJ9x1EWYC+TVlLMpGEQudhkK2
rwQKfTQMGXNMNUaBaSZa3qrP1LRYhtt9LO19lfZl6jpUv/AgfdsgGEJ2HoOwwiuGASOAYFi1ebIg
9nDfMry6M2vRQSbl9Z5i7EspTe+ERyETOwtR5sVpIT1hW31Uv2HLkwS5iIo4Ai4veH8LBapuyjNd
glQu5iSDPMvp/0rxNFHo1OnMYCOpm3/+b5I7shpPpQ97YIiDjpJm8+egs1Z8zEzJkSoRxF4+PYun
zCwvmcMBVUffXRpEi7YASGjFfWa3/WWnX2EkxDyERiX8J02u0tU5uU1Kg4V2uFVmi9Ca7P4ZyJ81
PRnDBj6ji3FUuHP9t4xezTi+g0AoDffXpRELYlBf8/lnfmV97439q3wc8F72/D8UnkD58gTtlOYO
HzKVm9TAR/wUrfmZwgWJuyyAvboBvMeICymU7VuYyR+ekZgnB0m/UfiV8IqGMHLwKT4GpcmVa1Mq
W5T/qukMASCfteoNUKgDaDsb/uZKuSsVO3mQ8HlvE6ldDRxqWxIWevRBm1Na5GUDfy9XQO7Sdbfa
kXiiPFWOqXtLUuPaNdCmmxSmzOWZS6+YlvuNNsJqvumhoNrDvyNITxBvlWnY1WAXr28RLEoH3RN8
d+Y/uhFB0sWHV9TpFy401U5NPL/bhGNqyH4bEkDJrNMkWjcT4aOUvljdtyQT9W4+UHsaOPVrrial
oJ8xQtuNj3gf8RpUuK9yTMyxM29pNFobPyWae3LkXIJLx2U4S97/H4SMDpBvhPzF6V9/wyNmk+8V
EUmucC9s4bi0/s+nbkyYbgb9fxDKdNqsEFg7euj1bGGbW3V86e35VQjZ0FRI6/ms1Au347W8jEqT
bIX/tKZoDdMsMnXm3lW4ehK0G3Z2xX0Peigerpc52PB8wr8h+M69H+UoUN49oebrZtmd1T5C7Th/
/WNOFnlukkd9Y/JbtcjGHYTvehmqg0cYHFZfrEp2of7goI0jJSszC6jFtWAo/C7PQs4KigKF6iFZ
bv1ApJgZgFqyMueZeGjBFcy2HXmH+m170wMRLWCjC7tkc4sBy1s/TbgHBFXmXHA65PP+wihHl7sl
IwKTU0bbiVWkOEvQwWhnNjlhIXgbe9kGfwwV9cxaUQYD37p2eOHbiZEdCKjg1eaTdO0aEKi/mTEN
Q64yl4+HZMW/WcdaSZP8vypMouxca6WjcASOfxkMc466aRAITi7gnHeUMotP/T7ahpbIZxrSPXVl
az0TOs3wlAl3GyhWUbWviVNCwcm7xUk1O7/t4Jfvx2QFbuvABp3Dp1AUuEvm7leYwh0IGoagXsP3
fSTQ3k20BzWT9eukebAlPPXEtIRvq1zSjM4saTj5j7RiAiisP8RQbd92DtwXXF8LOQ/orWBEXoW8
YAgDRblSGynDbITuy4woe9OorHet1teqrpTwyc2cnJMyXHLKEfqEaXT7mejtpTv/y0TVxA1FxIIA
L4pE0th7DZWzsBFa0GI01/qixmIS1TFmVwCLgCp10+k00jIDHLJjI7jj+mSybfzhOapwUTgpb6vd
Bh+EfrUiiQDynzz2vrGGICUof5tEehJ62YxxVXhtSdXJflRLrxRTB+RjOQaz0pC7ekF9/HYGmH98
RSBdafDhGET9DyZsAwuZKaoAF2ZBSUn4RA6zxXkNL8So5qTTZfwFbNqj9tFh8DHHyRLSkJtKylB2
zDYSYd9r/h2C3tbdEjsh+kfBfMgtvRReLcjYdsBX6THInMJtobvBN1nPgsii+Z63b5P3Xu9QSA1h
YmEF8LFgyhJ+2nHo52KnY3BJMO5qsMDUhhNbeAaH6+XXoYLNxbkvPzC0Vx9D2o/xXiDoSUN7f2sO
vypgHcGyeNEX9JdveneG7TgraUyOZCwYzeEwbpOTE9oM6clEcCn5mtOnTc2ez2uniWEeibs5I7bO
S5v1/b8FWYDcN27oqgc/684J/SO12R5A4qWvIPvh0iKGSjt+9A14uSfKVs2IewyR2vUT5d7M3O+6
piYlqrP6C3pi59sE2B06g0iwH/0dxf7kzSASXYssps8zPbA8oYdUl8t7+/E/HI3ua4+mZfhwQqfH
T8TWgVE4Mw73MXcZwgHvY9Iw3SC1U2bMrXbYiwyTgJ+4KSpMIzwawRr0HYestPDQZ3uKnMM8foja
m1m4PItsWMEI0AlLPnSmCCDb+FcUUaupZ8k19jIac/sEdyEShWfc1S4KP3JmC0w3lkTmF+7yYq9o
o+lZczvccLFw21uZxRd2cPJdQL+c62SUbv6Wa6+4yviJ0AOFKAG8uqNiK4NttXp0vg0BZUTMKddr
iMZHCuaKY3FG+wHtcLjFvEdKlxdjMuSUOno4gKo6/i/bndZnHztcHMHf/4ggOwmS914kB36OTKYh
gBbCfKU8PyaFvcHkAC1aiK7BxYVSBSA/1HmRFbo0cE2HpqD9do//00/mEmXHkNv/ZT1owYpBPdHD
yvqmGUAh1fVawtGXrdtNSqzZrvdZwt28dpXCj6UbMgJp9/rgtKqQmSIa8vAcpmjfT67sou8e3QmD
EIlCPSQb1TJz7FyY95rQsAZg9llMRGR7IPU3QO6lYnrlavCXD6p+p3LaGskwjSG/3IxT3kT2GCFW
chaY3VGgH8S5Z2dlvczvVYI485AeCQU/s2+cEDkjWHiwMjxPKAf3w2U90EyGeYM7ZYu18ZP5r5UI
HC+B3ydDjXg5xS/WAjMg1UmQafwzlHSQ7WD0j9typ2cGcyu/f/V9kV2pq26910c2Ut8h327wtOXe
eRBExP6BoR2+B4phGFiCVRGOne0NlSTluVWraCRYGSS1TQ0zXwZ6lrbzpNeQOd3Q6wRn7mx5YSge
E7IPI/XjQknSrmVCgUwQ7ffMe9n44i1y/mh82uyAYlq+6miKPqTg4ToPPfD6KeE/swJT0MVLeUZf
nqhXjn9vojNqL8/Njrku7j+HYa0xETLnGdHWNT1aC7DAf9josb6x5PKHpIYW2+G0JTWfebEe3oRc
BH+r5MlzD6xnSkxrE9negY41aOaQM2P2jIUSgLMZWFBPPpb6JGBC4C++27L2ohyWKJTtCcJvbZrw
VdUr5+XnDx2Zm6H2dGI7JMX3IUrnuhxwKgHTB9X/8mZ5lBf6ljq0o8tH/LI52efTymzLBk9andUW
7F/bge3afP64IlVuKnrdKIVPCj0QxkeEEimbVgOZ/ZbSYRrsiUrBaYPJpiy79xYkzRqct5jl5HsG
OZY3HjOa7QSgYtA8pJTHhtVuhd16J42yIxdU1ryHLJispAdyOSa7jKXaOZxZHE3SSgOvmOb/bcZb
Wku7QHGxaW/KjUXA/3wQ5lxC0Ip/2SPyE1H9f/g26q3Bt5CE7EeAVKoJoVEQWXpdf0xWVaW1iMTU
47yz/KG71XdZ0GjzwZN3CIPcrB8pfFmzoTD0lOmqoeypWzqm0hugR5mZrNDbgYIrebOxftEvMG0c
7CYVtLwWbEklWZYR8mciKV0QcjhukL2BCQ8+cDWGr30piBocUJlCAJ0sQzKFdqPy/DgaIJBwcyod
jm229tDD+/ldUwOcgxgzKRvu1TumFMNMUud7+JmOAnrChBqPeJpBi7lgRHEheZAY05Ym2BUnLGYD
+UON5aWjwNN9bqrN8wD0ULy4SMxvAhUIPGs1JodwCoxRDBhiFGv8shWhscZboWhQm9vYkoxNDpir
2IAh66hNbbSwqCYwh1V9svbLLIGsS7+H3Z2py0EkXl3/fLwjEtGzCMEeN+zR4txTIj+xSaw3r5Ut
tvgFOdsFmwhTgFt235zH2FLmca49Wn6msHOkuOJkQCRKshdG+N23R8VDg8srNde5rxfG4y4iz5WK
jgkinwEsI7cjDnxcVyFfk73ciIqX0uBYLudg97EyfNBXOqQoOUcY/BGVx3ilH8QGRolx5o8gZNWB
kX9FMsWetH0mrdS9DJC0pKofVtIZs3oxR4k5I6qgbCcpl2vX24fPxh3RNt8hI70EsM/CBM+sZnWg
mX+zc3wI45Ii+fe2YJd0BjZOo18uMVaDw+EvRSC2Ip5Q+OtgER7gflCWPvKdv/BjrOQNJb1mIUqm
1BKpmixdvlJwu0NXpb0FYmMFgCwmYMAJDJwSoA1igMyCjz7kbzlSrToiOs7Ng2qwvhoidoo84IES
gUdKuaJVyabWcVuYC5KkhudiJqlsKDj8F2hvLKDvB2lQ/Aueb6kKixxp0rQHXvtJ7IVSh3eS616R
oNXXEp1ZOlJ2HAU+VPx2NVu1ts54lCrHHpocUccVzYwpsj9w2tjIvPpVFKQyuG3do/fRNE2crsvY
A16NCc86a+Pco3XOd83DzbwH38rs39leXWnfP70ZklW+t5569JftoBZ8gcE2BKMjxGwXKmo/rpV6
KvfAWLC2aoHG/pCJSroklM1RXNTybIaHMBQ8X/GNmh7fOzYK5jtfEzI0j2sCN+otiebzb+Eiu14L
FfRMcRzUIxu8IcCs5mRe9qSy6RDta5svvKu26afHcSbcKiNNNQz8BdcM6MIGV3eRsPKbMbum3IvE
cSYckxseNTydXxEeelsBAonnKVyHGzM2pDbcSlmQQtxKz0gUpfHLTii+SbsDxBuTEH0m4oVtMmPG
xRyrJVz6qlx8nGsl7/PsevEe3rAjg0n15pyU4Cnf1+dWGyGUBaW7UfITAGr4V51agdJOLA8vFxea
Cteiih2b+vrxUXm+8OyFTpRUwUb/AnZoPhWsIBzzIMkMUR1U0IMsrGjYivBRUcM/lBJJqeZ0K8eB
WCX/4qCsttGwa4M+PxECpWGdnDRiu/dAXFvqdsFxn3NhjMlPAer3R9cZ+4Xvg91xdsQSZ2XUVy7s
UjAfYi00kQT40Xw7rCmxnGFgnFDmKOJ5oIMqMSG4DUwsxKqignvTdi9Kfx9KWLESU+q8DMynkdBc
owP1S63rrDL3nmoBrBwvNg1QGBu4AHjvu84l/NmXk3gjA/hukS6MxzHqcJWVmXVVM644toknd4nH
ySvHzAjYxRVqXTShGdc7DZzQPho04sWh5KhKw2ZYfiAARvCM0OlqcFDNh/E8uWaUW8w22vkwf6kw
DM4CITiScs82K1aq3P5Xm9TtbW9lVqJ3mw/ebMCbqCTqPodIIaMY7rOYsr/ivPNWDX2CsP3HTSJD
g0O9UQHPkqqAKigegD5oSnPW2u5Xqu41+IOZOdDuGGqQVfItrHUAqDp08FpHK9qh0CUB+F9UsnMZ
TLqLEJ1DVzPIHngsiuiKBIc1TdYD9SRRKK6ge7MFLtVt3hXuGLu3Qsnn6ZXm70cvO7EQnGE6/ylJ
0TouP3Dq5IzAX+cPMytVEhCqwoojP3p0ppK14crfd9sDKq1+eKPPMt+UkaPL+Ds6DTjxANFgI000
wsvxbGdN+qdsVIZqt4WEck/ShPmsdwH2hT9koPpFkDBPhD63x/KH0N4ZwB+A8b7nxPBdHPBwdfko
r1CRp/C3f+gANOHgalVk7AV5faoKoz9Gqx4JN53PqJiBfVSVmTayJJVQVP1hQB0rwmlXhVD0NiBW
ftohR5+aPd3a8/+vdOv5YydmG8fQSzCAENtTbdxdyBqfuWk3KRsPTGa8HiGsRd+hL2ByvQMYzAF2
Lri2yLZ1XXE8Fb9h8KShfRTPHtEeKLe9cRQOFf78tRqGwViIJwyQiN4nTwHFJecn0T9wayM1iNL5
M8J0+0QaevuTbMKQ6vD2gSYhzP/coMF5N1sZK696i4K3RM47HbU53M7PvyNNfxSJqrcUEBjBln1k
dGXKRn+eANi97N9MCd93OIHSNsmL21U34nW273KcuX3ah8tFfkzswcJfGWuMqbPvkfpKrWsNSDZr
2PFqzRpPRhkw/qopBchPqL+B3w8Fc8a7PUh2odqQ9mna0ZHNJZYs5+gTRNZ7yYWQQMsW1+sAKsw+
w2PnYvMAdTR77YydVY5ma2XJ8FgQBeszq3qtPccnotPnYqZcZRM/kw+VK7PNJgRPp6R3cL9y7gYu
9YgRVG3rYr1DS+IXmInLQ74Af+l1yow06vu1zxEZEGudw4NllMnw633eAt3GNTLZZpnRIqv0llrR
EClIc++fxXrT0wgXThPVhGk7PGv7uJj7EsbnSWbHeFCIrKbv3wYYFRykqfjXFkr5RvwIgD7C+qQF
ljy9uA7yiWlHlS2j8sI+SWDaWp2gcjJWmJ9cMsTxt1U5ZMcTvmHQRjvKVu/cG94qQk8tkqlUxfBk
EMhbbrHdwVTSIo3ZrcKghV8eok8+bUu/1vmLfU6VM2in3hItWwlN8CXS4zIwowPTH/+A84EjrWIE
lRMBF9xLRAivpsHKLf7GgipJULq9CCBJCiTJGFUwxZ4gDoDmfqHQn9IJYNCEh17brzMVL+uKguyN
veCC0u8xPRjR839eUjnnnxOZIiruJH3zpTkmaDr0XaIdtpHUtLilmkrvzrf7s2xGunPljHLjmeb+
4AyWCIO7yeMWfG9r/EO8fWJK5qb6qZCfx0w+T6fbp8y+kE7Iz4W2bK2hGz9z9IjdEffHMdpTkKUa
fP1jVbe7Quy+r89ZHYyUjQMCytx8UuhVTalAMnvU9FYmiagkpjU1iv7vtOFGLrYOqtCzXk01tS0b
6lqQgOfACbDMPQg9lOXCbYSCwvqcJlI3OQFytCkuSXAwK0NNoFCgV+NqWKlJFQwKu08sjmaQHO6x
0HbaGKBi04BwqqOqRThqieE5nm00Nwk/artLzCbwDGwUf8CiP4J8n5ueeEDFYLwyyjULEaMZ3KyQ
0D5Os/u+q938WAgJtND/3fuVBdlaQ9bXNYlBdQZm0dupCbo4tUKyQHwgc1tj6xGRo+agsvNB2lej
RiVJlmtPI6wXZtk2W6/Qy7iuUxPQrwYa3ZfOn4v14YDFRiZLJg8dztvQRIxzDy3+R0q2z+Ay6h//
hQFTGWHwMUFD7VnHpFOWBwl+MZhi3KsoGmq5L9Ha2zCPTQ0wCpTkFpoZqCIhDEA63spcO+UyTW/2
D5wIYjr7GfpH+gCFQNfiv3jaP7Ry5PTUoRJWdGwJa0n6uQIXP82AkUVp8SQ6bWX+N+27jBVVmEDI
Fm7Tv5f47UvNkUHKhaUapSN7v6xN/5PYbWXXj1LDKoqGm6YTzrip3YXHXSmSq0a2Yzh2IFpGBn1O
GiieSWCadWpFWwmhvB0LlijCmoLOjJmcdIXv4buF9bHwtdGJ0nEyCybf9wnss6fwTlA8CMAWEmq5
7pu+dfcAXMtM4WSanEdvtNwEID7ibF8nGO9JXvTtZNPxkOYWX5W9c+NuO7IwsVQoG4CNgBci/CmI
652brVfawqCvcmZdVW6ngn5mFEtV/3v00blD1oHfByoe4YJ6hWcoaNbnkjlCEqU1dyRVYDSOnasE
BorV3HHxUdXKkFrUTVwuVRwxwkLKWfY/69FZtazEBQcDqznDGhfntO1vTLfHWqVZqdGBY3TwmpVZ
hi0de4cmndb1NLmEisJOOKwZo/sNT7qECg2kFMoQjJsZYjPf89xOhfaydeo19KEqXEosOZnAI/ar
IzMsRnfaf7ZrHIWrVp3dwYnfeBk8snP60ml5bcqVpY1tYtuWVag8HdMDtDAlgMqHfTk9he/u/r57
qg20MhWfqokTAwIrcAnYA5m8n6XpvQvcrURTkYUEpWGRhz7/ECR53nJhj3IhNQ5pfHUTqZBCtsvY
+8wj3ZHHXnusns4SJMeGkESkuK2suLuxJ5mSaQhy+RQy6xtwJmduQMnXUc1WgzNjCLHrFaMd0f0M
zJgVOt9nXE5n+g0UHvZi6RrWFrinzdEIuLEEnMJe+Q6j0EGwwkwY3k4Wd0YTWIcyMYrXcKlLsVNT
FFMV+0d03i2145lcnqLPuQ+dwBW5gXEtjBo9WWGvf0gl9VRddfEjeha7V1O+vaWZkTM9uUAq+cDw
5Bt9HSSUUrdTQ2GJB0knFhDVPole77m8MXTBilpD1IFqaZrhw0QWxZdhGz4jN1Rd6pVpN2oybcRT
uT25GWwlxJDP+SefZwCT7XUiQt1LHQqvPayZAUrwZJ+mWcQY5EYb8Xck6fNQhyEX3zJzWhOp/qg5
15i//fI3ueXvF27EsZ5lbKPX3GoQXLQHlJ4yfrJ6lC5wJR8oUEZ5wun4Y3t8P1p7CYXAeLUSW1EL
arfmXH+o/fvOfSjQDRXjuwL/bqfgKOmDqpziJ2BYNOBAXImgI3F8bvFLRnQ91lJ+CKoLyuF8cWA6
1oKMdYEzWZaHeDI/W632cHisqPubby56UTBpXjAmg4shFNulfAcxRTfJFF/BjCMMVT50sh1Nd7lz
GzNao0H9TjPlbEADq/jEP8cg7nD8yufPLptzlUXUXg44MwtRRf4YO12bSNCFet8bNPEVK+xmzrnr
QmA7ensZS2ktbYS1tTIo3s+y7c2Q4pVQvxvmptT4fzONcK7IabPWgF2r5sbGZRXF66U9UI7ausFs
TOdbhQNs4DH4fXj2IUaSRGy8qQZV3okKLmWCRboKJW7ASdHpGECBG2G5wV2wodmbjLPm08fEWeAw
+RFiIyCa1pWpdiEBeee3Wf/V7FNLJllUYZ4miLH3m5nWWuHKV2o9SW2U4EEdkJgmYvBAbE9yJUAg
h/WxVSGfhdTAbB2Ez6mRkgPdaU5Hv4Lm8sH82USgD15M1RaTkTxwZgNMFdAxFadxAOYhVBr0i2De
mW+NGuIy72c4EY32N0uBrbbaUNhEvS0r8KGF4+HdIRFhpmgGcjVNxFarLgBDwRv+0dlbFaj2iGWU
0TV15RKqrjQRSJCUJAweIchfD98chflCZNDeOSNNjm00ZZpRKV/c41JV66BFb/FnnQ8D4jrytkq4
CfPHQgTRy8i7PuSaF26bGKKBH+iRnoWvj1RmFqg6NUfT5eQSH5lD+u3HSDU4aRJ/EgJc+NEoaMca
iEJRRKMReLu2Z78H0itpUZ+vF7fln/HUWM2qTR3tcnk9y6rh1d5g4bjk7KWFvt1jHILfxqK65Cht
Y5w6SCDheV9pBOHkiOs1PA7cH6yP1OXg0iUD+FHINyn3LuSdpTiQLXEj7rAeiLCls8MHcsfYVDVV
ItWSopvZ/Ouja43VYtctZXR+FLsVannP1nCUaao1EN+zpEA733Rrw/SlzeUn0tb8wLam7f8iWpN3
tArXVNYzrpZtI+wcpVVpeewaM10ql+llzFq8WULF86ssPdPCsvdVOIPzcPhyXC8f5ph7BC6jIImN
sMoD3hA2xUeDmy+n8L+ZyCWiMlGjr9OJXFCHJJP8eEHs7v8BObWDtQHxQoL9UkwFMJwx5Dh9SI+f
igIeaGBDdzWbdN6no/vgOXGRkccuAhwEyhKCJd+pxYsEn+CQgCTXgnavqEWZArcEo6s+NNXOGacy
oonPJq/UvVeJDVVwKTENHqOuYF/FDa9/yKbvPN1Volh7LMrideEHYXsuGydNj91+LDrr+kBt1QVr
vUqpvqZsG0Fe7xu32hnShPrDw0raMGGCHyDmLSOnxVu6Ve9ZD+BdcHMN1ied4t+YOxMU36b3seeQ
97qpSeThDZYCMBttsGYejgET95BdxP2WzoXAfISY7oiRL46UK6Z+titfKKvGLXtOAQlYgUSlmiNd
Y9tFoY1h9HiVFbysv6yxM9rx3dBkOypJhqvFV65hc8xidBZR+e6frRyiCHc5cw088vPNJafx7aPG
WqdiirrtDrFO/89JUWxg1aYIeNTyOSprU17yWZIu+bvWN6B7AUYfu11Fvtz8j7wZDlAD7YLL88LX
EZbc6nRtSnjGYWY0IgLyYbxj3e0T8jovKxFLKv3N+nzwAztu/GyJ5yTFl0c4r4zhGMH4/ANhH+8u
NL1sWl+CjfmRINjI6z+J03/0AVeJ7ebKo1EsTgoKWj80ZkCKLo+8v2d0aZTipuVjxnJzSGH+3AcW
p1JvNNCSH6YE/7sDK10lW7dGEhiEKvcKr5fduWT+S765WMido2X2Tg9N6ii36Q2SE/Zf4xvVX16D
sozi0wNfWXK2TPBtoDNxWSPZ7rhSQdvshXUELXHMGWGTqe2LEBzZ6zHv/LQ2qDCEZsWltzzjbMfs
T2ajN8HAnKs3CUrUR7NqMLSu0bEIilMSQvh9d+HFMDFXvcYnMarAoSm3ZGq3rpRufH9chzxZ60eA
9dv9cfeuIeaS4r6NF7LA+qu3Sm9Hnskex7Qc/ts2OqeFoKOsl9o9q7nc0vWxwlNo+d1EhqXnGQwB
D6E4TRT1Y8F5Fgou0TNp5a8ugBZz425uzqsFRu+l25/FsGntWB89yieQeWmqUDITpIg1Ma0s/yJL
0B7nPhi+34SHKOi5R/pt7OlLJxLf2aaNTACjM3bRdxzrcfYPcwyUxsvci+EMpk362Lg70nfFStU+
leZUCzNyPzmIa33UtaKnQm1zDOw4Q3oQbm8qAQXBhq9aDQKHR2lnX+qSU2xpiCyqWDoNoZDliTdw
92U6sCkXN0hWWfa3fKSP9VaT6PVQG77/sR+bhgixFNgtaKeqdYPf77mw50xf2vhcxWwXHrDqGf3q
ERbatEucWwow4H/XBUEBKJ7EIfz2b3gQcu9/mzYqDKFcuI5TbeSXx4x6YdywOpEuPKgB8PBS4q58
f5RCyW9rUtMfQMbBwsNkQt5OFBlsBW/BFIBocmnWFHohhkGRbhi7/SPzemAAOoHHmXyjBDCh24pG
Srrlj4DXNK3evkkScSiuDPl8AYpqoYJS0arXPXjzEDzV9cKNOlPvzVa7lZVOGULNCDFdNbvcVNtZ
Dwg3Gl4QQEKBYMJfPx0qLhoZ7eFBp4HoqrIqsIUu44aKqIf5kjlQLEXWl+Rp1RZJcIfX1RmPz8zA
b14hBJBliguZQqaG1OI7uy4xSm6KeTEisXyM2NBKrxkr/GVqdRtD1Es0GXOphrPYGIb82l554NXA
sX/c67hogqG+3Ox/v/BfifmUCvoZhtMgd12AjwxU5qNO0LG+dY152M9GGf6jeoZdrAk2rHAUBuOR
vkCgZ5lBS6lB8cPt/bOHR6836dc/mK4cWOt3yQgz61WXZzUfpfpv7UD50mlZjNcI0OHBSyuXCZD3
QvWNad3JEYsBMA2aQerR84ZuvETvL/gCWAiLI3ehuz1c4Jp6efaBy6CO4HmmVc80zC4v3cSSmLZm
Vd1cid+CRgQNjsH+0qrACGXzFeUvVT3kUhKQeWw2ByfvdDRxGbJLpXSBOxLSx/YQfOTS0FoeTkYJ
6AgSvGIXBvL3qvdBzJHWAbfey2NI7oTFE0hPI0xoB19usU5PWvIDUduRSneBljqHOpntyZ+CqV5V
MEEHllFv5quZVSKmk0MaKz86ZWUuTXGmPKU4ZVUv50YHzgRll5LzLjKx0OiXfH8BwUkONDgXSs61
RdYAkGPP/9oFbM2yAHBHj7D1dOmXr8GMaPv+mR3gSm/497srt0U2CAqydiYs54rBcoxTTQ7ptwNS
+upuuxV0SduBr7xA3dx842bWTgU2s8cuXJ44ULC9Y/FIr86h4O7PN6ZoQwgnyIWJvdSkq8eOBdke
OeySTOi1M2P9+/90VQnTXywg0oe0UysxUIhnaGNdYfdMH16yjhmBbqsE1u39gnH6iyr3yOsOTHyZ
L5mvv9ZL+aPmWyl/zbnw2QlwU8b5Yr9dxlXBnTaCpH4cm284frdapmhoPnicLDz//dDA/XFyfdNA
qd7dNSjKe48cZmF3FZmLAQSIf667G/j8yrBaKGHltjUG8EEO8FGCrrxQ28prG+26MDIcww/6hhTh
gQnhd6XiWvwOW6fVmA+fwpq4TWpY2RseAsvciZjU8/2ziHYjH6vZ8Qwzi0vg48FOOJMmDIyVyHZj
AbHSt0I+F9SFRGjBK+GzO0Y3HZnfiwtdUzqAxL+elrJ9hHuY/xSV8nB2mqpKGVMwAp/hYqcAcTwT
JJSyY+pyZt4C5LUAVjh9duQwr/ZWjr5+ZvxH9NCJ3ISySXTv2/WhKiOJqJAEhYDpQWmCyQnGFdxQ
rzqlTMD0AJJ0ZgPeQ2HD5YfEyGfqX98i2qgURpu1o+NyrnT9IQGVridHZPiPueuZT139VzbbwOdV
GMgXLTVs8JHwz7GSiAcjRy5KRPYvoadefc7Co+C/2bGEjTUfF6BivrPHAVfjaFismZGMxdqS5Vch
6yhrlzkMWhgt2UnevcwFceXgE5/STD8nKWnfqMLzJwIQIySajPRsg8ZO/cq/RJgBTw5DoSPwYa44
8ZWYsL5WVAQPaeHNdGdZh9D3c/8fHOiT9RLmtcsqgxcooapW5AsZSPrXPCgg24ZFQq/GhNswRDEL
gTzUK5c/ULnpMZCornxgwum4c2NFLPC5k+wLpVFBwmcJPNvd2ADphEMENpn4YTiqfR7nSHBOkYwN
fXc7oJUtK3rNc+v2pLBzKVjGfKSSG9N2CGT1OyXVXbV8JJ3ZR2BWIeTO9lmaygMBeHBW3NVo+wWk
ALXOe0vFREu0aPkUWdqV8KlyPHNA/xtx6dzy5T5vRxZt2dHdERc0Qgs49yiHI7C1LS//t23rUBi7
KxV07vEMiR60xRp15QaBe58KvLDW7ipKUvTZfGC9BKyaMCMH+9WuMJkMa/BC1okV9B+yfxaCnzEa
1Q9RRTdWc90lxaoFTe3DfGhmjfb+lF1nIm5lIzJGChWGp/TlK0QkXMA6V2fUwvvjiwjmHHzd0aOk
Cn6k1iIz/wNrSV++m8IyVMK9CQWY9ybhGM/2AjBnfQ/kJea38VmWhaC8/kv90brPvR1E55mncrno
mI1jk0oQd2JmNQaIM/ML/bKBJhDsI0JC6x4CWNl8UPZ037/XnS1+9m1ABkYZNSBgBrD4zZpYJg32
qZZtpswUZ5S/KPMXduVlxTr4aNc8Mc6B9HZ2Yq99Potoa7s65Ds1BPFIFOGSsUlCar5hGcxdZeG9
CzKiK5WOa8ptZRFMXeV6l/MMKJFOU7d8RSitTXhbZkH+vwmg/GuLOmEebtphhuq6L5ZC2bh9dF4O
n/FoyHj0kFWkhPZhjKpa9mxvIBjZQCGmR40L38uh3jO+SaY3Xct3AuTVOuRrq4r/jduaJmKEhSWg
UpNrE755S3andGRVBWcmV4MMcu0lgvJZ2ksmVKVZRSxcsohQezw83xijFVuOF22WuFO1yEjElM59
ZxlITo3nFdeTAMQqBm1ZS8YFdFqyuQluOwcH49hrv9ePGikU9gNN80K2scT1c+PIWW6NVJr9mQ2i
mYVKIVtGV2pdyRRtE35q3w+/fMyKNaY/osRRetj4YuA/zzUvW1zbg+Ij0RJkZuDO+TeKtXlxAsFI
z86g7CS4m5uBxYIexLoPs+zNcP2n49LuPOCqe1ncdwuXR8Dr35He/pp9s5Xh7N7qSE5Yp15dNKXE
cmleR+47eu209VxG8Ae15YumLulRQwZXl/tdmc3jVz7D0V1wIv/NljHtRJVFTJ/MphEpDBweew39
PoLniSqolWQeF3aMehXgZqyhQOds/GZqia/6Zi999wjh1dIxmbuacdeeHK8Jzkx1+sA1UmKjChhA
MjcINFx58ZBhEzRA/7oV3SqAe3oymAepQXLPe5v7mIF0q9iMBFie0suLYGwowD0XqG2syT9Z9m9Q
OkJez2UZAPvHl4NjqvU8pe24qf9pwWVNqLuS2Tu5fdnZFCsi/Iqfp72e0G4r1nfCFw703SA8NYRO
7JUGh4T0H+SzAKSTxiL4V+oXahoyr6mgq+YulQ9voKl9RMCcQu/JU4Wtu9LCqVxvyWJ08lrBCQq9
jx5DvZ5NnGh3PX1iLVczLtS2hErSCpJa1M3nHFhClC0VTEjPx7akKupEabvebSPE4Sf5D4b+aAwg
Q8APZyTit3u7oOS8EAnMmxq7EJpoJwXDrrInMAF95v2knk8jyT+Rk862l/xM+Img6bxgCnIuU/0B
Vdz2KDhks1K4K+K1u1+k6f6t2+LPqrbN6BuzGUPIEN/aG/pbMzWL2Hyl7+wWsGPSKefH2qqgeXDW
+19/VyTex98bp+G6f0KEQvet/9+Bpu6h349phS+MVyxrbmo/UX/elNC/ScP8TtcEkuCaH35XpVGZ
FeerlmQCTfuLZutwb5UABtQ5P21KYuAA6u7gRgHi0i2yDa9oNYhFvcztn10iBP07LixNKefZpLZg
FpRYM6/Fah4SutATaa9VT1c1kSifGG/oTih25JpbV/a9F4t9Fte0Pu+SX8t4woyNOPxqTnPwixK6
HpPZTlv7CoNriSheRShz0ZprD5NEWPaVsNv2kOzgOnw2j7lzbClClKV3RxrDlZ3Xu9CEkKOMNhPu
gjvejpwCqdy8uRPZUc1M2PgJ8BdyjMihil7l3g27A0RjKE2QHuXVqh8jwV2hyKbE/a36PM9ynJTW
W9va4/E743jykLdVUGEsWOsbeM42tD9qZBmSyr1l/D20jHHzpHtoni+EfUIfiLNcaWE0PhYaVKiK
Y7k2HbsH+uwXdKa+QkhpdysQlHk9nZpJuH935uDFhJvFMsW76yTuLhcXLlLOpn27WeAsYQk9Hpko
UkgnT2TVgoo8G0ajXBuxBnFNv+KybtxZ6uJEZRPbGS2R03sNR1owYwwLzZHBSw2LnAgrZfCvo1fk
7jI5uLX8EW/X9+TlznlwY07QQKP/w2La7/iH3XXtRsdDyN6UYuQnKCCPx/Kj09Ki8XRJ7c9b2Yw1
MPyjFIE4Vg/O72rLBJHuwTs2rx1TVj6id9x2eJnlI6J9IWyZewNybGG8Yrq5VPcorJgTyv1I9hxU
yvL2o1X1zcj3p1crv27dnRx3JWfJreCwf2aOXcMonZ5WiulWIyPVOAYml2TFZXGX/w3gFZ1U3dB1
nCkVAg7DTKfctX/2bjHEsGJa3L4ZLwhI+D4N2o4k9feue/Cxf7G3153jXiAMbU35213QYH6plKNI
FBYR4V5jVYUrfuzOqfP7IkAhdBphUgoTjaNVDmrk24dHkA7wqWMypCtqBvQ0ojtZ/VvPvM7YY07E
5SbhNRvaZOitEjRomz/UVeKd9njrGuHIW6GcLM3wJEKsPSwBjx8gjf7HY1+a6mM5PMqH/BNcWOUP
6zPIHJqRDAT54G5LFlWT75RcqDDAqgJCz1+7Cx48ejxovxAWHHqBp+2ek39a3SagCNgriAyvGUaH
UeyTWiP0LZ7B1K7Oi/iHeur0cgWW7yKHyaFMd24Lr+UvyGcD3qr1ujnvxM4OGjUIXKQbQ+qUTfoM
m2JAHdWyzyaVNxleVw2y3gNO9eS0NhgNc4Fb10koy4KLYKQB+YwhI3bgKZ8ic1ME1R6RbCzL+nkH
3rKYLjiqxj2k04eMJZAcbBbam2pLrxDx8ogIj0bj++uB0prVJ/stMFQPNFhOUBMuDGJ+yDn1tz57
v/1WIP0NBjUSfdnkVGyjceYrVBAAb3E30PKbmQxbYIvXjk88YHRgC/+bj1DXeb/ABSEH2/ThJ8ik
75fRqpA+3ZUzk+PZ/4/3Q3h1GliUkiTA8+EsDti2AefkBw+X6NSJfEU66kY94nmvTYuCgtMsC7r4
1azGsCwDUL/iqi6T0Os5junApnJVGPraVShfYHvmGC59zX9rFQERsTyfpmoun1AmTf3Eh+Gc+C7d
IgwHv27p42I7FQ47j6MANVZhV1HOoj3VdVAuJRDRhCXxY61CB2G2PNdzgF0a2/izI0old2J+qUuk
KDvfjhzEbdYPrDA18BDOxdSSd0PGodd3Rrz4fNztHuBx29+UO1+eZ2c7rhPwB9JaVhhE6A6N9E5j
SC+g8zTR1imCRSx3fHDYAtWa76M/PNDWL3C/mkGs3Dju2vAGARODehQhAvnzUBTJv4M6H7Kq2Bvw
tsbox35IeP+yxkh5NDpHsjgsO5Ps/g3tcP40Owpe2kaZ3qVwHJaZh4ASp7pHlAvCUzOwBwWh7cRa
WRAM0aKt3Fmjj1D9/H0tyYlgWFHNciOknFXaaOSCofzsN/dtyDuV9tMc1/QzAisa/cirbuvk7sYH
kzORQrhR2lfkEwPIy3c884ZojCsZt6lfF1uUJ53rlT+Q0CL5wgksQeyRoUIJ14V6nkgTda/A0AEl
Tzb/gVhAwnKNJdxHVBKpqTsAl33jD8Gnl3oPMi2W/okC3A1iXXWBD3nSr/ozdyS5G/SzMgOF/w6Z
o3H63J/L9bctg7GtCaq3k2mbyFNkWYEGBcOuPGDl55IcD/U0aN11kaoV3y9eeMy85HRbWd+zqXCS
re84jgC5I1fYDLcjKeQCnFWoY/8T2Mgi3Em2MiUWBv8yTgHpgWBQXggiBJYLqgdjbg1FXjL3/J+r
ehEWRuL3MreNJWxR/uIsF7HUVTSw0AEG5vpwqGhcBCVJ27pqGb+BznJHyKYqo8uI6nXQo3ZHYloB
3IxwRnQKGfkaEKAmnkcVqyDHXeLVmByrHZORQCegxNR/Ng2xeup2dOO7b/AZFXHnm+izFDTszk6o
ycyG/McKb3LUKc9h+6PWj9+l7eHjw0SRi1U02wHhoeHzohSIYAijrJWnCEoQXsLA8dhcVQQknaFF
GrCnBOPWB7/VCvp/MEdy0csnyn2TQTO+JI6dQPXxesvU7fducpl1feDsGWozx4iE5HuxmI2JCWG2
zgm6FHv4VSwUKpIGp13mtuv6gW0uUG30AADs/Khi5QhjMF3kOlRWfHDie75B7a1fXkgtlODBD2Aw
W2L7N2wrYia3+22TVFSG1RFIyIpEaYBKAZNAx6M3HCG5Ee2GBHKBfwH7bPjiTgNlmhT0R3yOx29g
DvFfHiE5WCRvg0kUoC2k76uE9MoQigFYGdxylfzTf5+99In04gVvTqdBNc6pe0NUSoXlLS+3O3Mi
MIhreynsaQix+gc8laa1VquxWWPbT6HV2r7eIOqvE+4E6V0CzNYlgf3nCKbrLN+8qjynj7KTmu8e
mEM90wspqPEcqIcsxxf/IOZiKUCLmOGYwtDRC99A2CxaIUVpo4y8ww+Pv4IGEhkjUOhqx3nzXe2o
/FoO19UYmFFMUiEComngJb3v1Xx/F/IufEwlQMAzPhjMfrvXK6xVfW5D2n0TuWsCVZNIH6RBUhs7
PW/6LpHKmDpnOghl87Ch9BU1SOH6X/gp4svn7rDRJbz4Ioa/A2pNd1qxlgAJ0dqW7tfSsVbKfB29
yqUzgChBaYjZxB2f4afFvzQFx8HgNFO4EHVMwcCGmbT5KlTfZXhXRLIDcT3ncK7QiO7meV2mCM+g
94x1YidYNB1P69vCtdiL2Eae9TpDXKsieUqwhw363p2YeMrlGRWSeOvPmpUnNtUORdR6N/zdrIPn
mcWjWl1AgyhClpCnwTXTpBLYESAJNnLaONpbW/t0WSIhW2BbT7nUoBPbGgDr480Mm57mS/RqrbXT
oU5WSr1E0gmIZ4xr76iRG39rmoNSaOsB+rtmvHd0Opk4rmolqpsJt78pfHNO6nIf4onOhE4RjxBj
jRmz4AhUr3aHRFiri0bjX86w3CKL38SHmgZAH5VTBuomHrJlmcC57Fd/cLST+C4xZmz9aPjLt79/
nQoQx1tve7jSV5TksurAHdd9OvG3fdOffox6poHAvBIRpILUnwkJnirElgoJLboCC6YDl9ANKhWr
G2APFdbkaqbc83HdzqgzzT1HcbLZTUMcHjfVDNJEcIj3hxjWaU1brdovyYg4ALGkVhnK1YJHM1SH
4UnCSGj/6iy7zqDPo8+2ZoFKnj9f0PnMQiNMwA8tX4Dvh4HJLY9PCWs/Z3uQkaaTvhSsVYFOdpQV
EEPHVFtVOg3wR05Uhpoh/f6Qm7A7sIGVvb2vPIM0s04qDOM+6T/1By8UwIl1oqmzhWpNeXFxAm2S
MQCEF9RidToKhXRybjHHdViwKfSb+zTdMF3a0Klhka+bwZsnYheOxN0bxtZN8vpcNXchg+lOfo/E
9NdUgkiC3lBlGvEpK3VBtnwaqG2tgy69OUMHYvqY5HW/YHjJE4+Q7TZuPt1G2Qq89OptFMU+unYZ
te/Q3sPRZJ93cZDNeO2zPdy/gtl3ppRKay28PvCLVrPlYv4CJE2aHGbdfAtlmIAmztBcg0jciwa7
d3wo678/I1FEw0+QuEUIl0iyMYrMQt0V92YeaAyq25YdLm3J8mdHwAbiS8o458/wB6Yi1f3VSgY2
IJ5B/1bT0vAceRks8aIixFK07nKhCHr8ixml8VpfwyZIH8Y9NJGYOy2nAi4dQUWeWr+iNl4SHQ4+
K+tSRBO4uIADcCo5O/+Tuuxq8he+1BqsxX6zPTzVzyxi8bM6n6nzUNsa8ebOvwgmdtu13Mr0SNG8
2tn0V92SAK4q1rBHgdH0tCqubKV32uI5HxodMaItVeCTheR+zLlsKjO/dfDMkSNaiqFbR6/DwU2W
98b7cTX6rJEWfy750Un90alla1Lc9WyGnpBpmUvnB50DHLnYED97GAwF2/rjM7bnJJh/qJ9xhX8X
k3MtWz1aXT1Yi4FoqBQ7ACn9juSqiJ95DvTFxKim/xSDN1+9ZzV+2SSn3OzRyGz7WGaCztRFCGnx
pxaqMv5IWPZm2DdevJiSdYOPMAjZn3suwpCD4uRcTJxFucRarjo/h+jYn60VZWZvslkaPLfLEcgZ
q8ZGGEalHalBNWTjkLJ6YQXaqSfYQwheFgO4C6cD5zaZvgBDaBPuIV8NJStvFy/4f6I2DkFsu8Wu
N8YItp3DXciZBHvkh7ZxoNX1u9JnCyucis8Xa4b/hxKHDM8EHLtW2D75dotsJDDF4JjAd4wmFSq6
WtrIJogkVdXSyWZ+5ep2auDFPVWItSzNY1gvkl9s8rbT2ddBQHh9F29dAoUJA7Hl332HM4tH2k3a
ll8kxRDVEa2wDXH2v/UVIOhHaP72AUCVZJDWwx3m0VQk1sW7SmW6h3goLy5yLIIKRh6clQIt2Wlh
ty66e/C7Khj11U5ipBLbexWslrMCLJcY1ClyoEA72hxbXPN0NZkw8RAjKNFHCwIbKlLGNBd/Vrsh
gm9jgJC94HLkWgMeWv/UzNmiqdJNTbNeOkyDeTwcv5IWNIpMxzQBUcZa2F3jVtBqQSut6ZqBGkb0
VRTtsjKmF6ORZqrSYbo12bgDnsFsk2c+QkDYStXT9Nm5INHPoNkWAhgiEq2HDokzeFqXkrQxRBuK
J3DseaJy9uKCbn97gRzGP/DIQUulaQWTvDiCeFl2aEuEMisDjoVoNbYnYAAv6cPZOUxLK6INWzkJ
AevpG61RPWukqyfUjO+qnujX0VMW7bGJLmuR98i7yD39d6sq/tjbCFy3QBZBxNlwfnP8fUPpNyyE
9pGCLh7ksB/i7z0cR97rcK4pNDZ36ff2Y1gpwN0i03qcxdevU5N+rk7PgVihGm/ntg+9yu/Kupxj
GbxC3qBd/CeLDO7yqVCkKxPIXz43wL+vyHvr7nefxhevDDHZdSm4stlh8azEdWJKYA78sMlkGgTm
CDQOsAAKPttzTympj58H0VjQ2Y33tR1yIc3PvdUbgmBHeXnTk+GFgYkgDDD96luhl5l6/Nazr+mp
oKULz+2lVG0fytes5UbY3VzkwDIwGkjTrAPa86AAcp4cze+jww+EoURXA6ZzzEwDkaF50BrhKnG/
swczj0bBZZaUIeaMFrG48Fm5UwJAewSSPiJOquyiuMyfEICDF5eov+6bi93dZvU0v+NMe35n5W1d
cBi4Dl13U0/rL2sND7dB6PaccUvxeblkdRswREthl1hZUO4pQ4cCL1Y9JLf+8pLZSguJmu4cLk4b
1hzDa0QRQ6tR0BTjHEX9T2ul5fBJlxWrhSmA5NGFTaN5lmrtKrX5fNcVTXIQ9kyMPXQ6AK4dCIDc
gjAh0ZLN5qnnN9qgIo/DG0aEZs1SL57tj+MqwijCMK9YDxxQRglztWfC+matJQa+xsveUwnHhOaJ
LCH/F0lWE6AdmbukHshBlRMwDzNcHDwlCw3S0U/HT85I8ih4EIQ+d2RMYvUjYAAPGqWS7KnAEAh0
BD8fLCKOROrpxicIGlKPdHaAb6NebqHW9gEh3ogeyLdcgrrW3fnWct6LfA++aXx2jdIdqs15T2v3
Uh9z+35o04KgoWtqnDHNO11DVXKQRhYxdEweYNMmSGtr5kfhGtGcKTZ2yhV01Rp0kuOy8XozzRjh
FGPGak0vQfZHWTRAvmHHBnd4d7M7PWDgZw0Adh7aLyDec9sHml5KCJpx4C83qWJmOiOWp8oEq+rg
fwG0e2TjQPR5JkhRrfBror3lZ+lWhao5O+D+PzbX0zodUvfUeRyOfJzYOwVzIkmIfJwVLPjVaXm4
HiXV46X/O9HRNn0Qka5YqeSu77P8Raou2dhhlWrLNkZ7Y6GTS0Psp2dFdGHYC30HcnGh6gk/SK48
VUtg9qMfepZKadykr302I0a63WFSw7W6H87Cg65y3d/ZbotRspMKEQdPfGMbwKXgE1Ru2HCxHZVA
zCQ8kOgpPEUpd1/+pjLYUFGjLHRjuJ93httzVOrnKUm12fjaGjqKmwJE0n8EdZNslscxzVwUlfoy
TnZfznn1/Fr8B9ryGRELs0WIFovyDHK8nT3eqhXjUQOhd5Mvd5/c1uS0Bhqc5ehyL56+NkZe6e8t
C/oE2o4Un93Rjzp13B+Q8xz7B2VZKXkvVhh0vahjgBcRVyraYYBvnRcUP3Nf1B36GoLP2q0JIV1Z
IDYof++qPrizS2apuoIzPXKuQM/yS4M3WCeqyKFuJg6vXQDf/jpMVfoxXPksU7cQMHEVNxNtMZys
z/Ad7luG3Z/dXPw9B5b8ffKiJ3nOjusSZIfBktw2Bm/e48ZkVcl/oYtoYvGGOu1fwoqorLZNnJ2N
FofjE3HCNFYUG2D2VyPA4tJOaPXTqIAqu3pT7tApA7Mj7OireI6ovYx67+3PTi7Ghp2YI5g1oV4a
D3anDMmNAZ3bSXc4WiIBlDtAR10YhZhyngvcb/MwTu+tCLcPqnOB6cXgxLKSokag02c7Uh3jAEiu
q8GEyhBvl0LFjkUfEdRVMggUr0WaU6r1+3zPKkmQDh516lQmkXF010y3gbjRf8oloXp9dryyM7h4
2mhcOlwl9D0qOodwoPFiVd8Bx4ueleph/QX3lP9a6177Q4nfxBJOYn/R9G7bCwMDICzkoLPaNSEM
KxT+nDpwnTV/XJFJIBrbbbOLPyS8dIHIq6tY6v1mAop7DZIpGrf97bRtCES20qpCyRwLZyDCWByF
74Lym7/uom+qLsDJkU1R1jDGdQXYEkxvzblBUpaYTz32KEx8FilZNzyj9+DAl67Ws+McsGkT5G/x
zD2JopvSxbZjw3zaDtNfRokQtFYmoo0Ag2KhbDMIIQ9Y0wN0iiuOxkn5EFuMYp/5Lth/BK6/cl2H
EjOW8eacKuwFDVe0y2aLv0AknqqY8Im3DvcTxw4ulG9plQ0Lp/oE0j248uf/+0qwnwor/k4R5qH7
rL3lmY09IeoHlZL32PQOXmFdZ/CRpGQ+VmC4RhIBE0SxS+3sCgIuPQOWhT6NQLvcrV56CM5j3z3i
HDVwJ2wSTRUr5kLxSkgBglIDrhNlrZ+vshvY2prJq3wk9On3W6nnghSoKc5WRIYu7+uC3+QAL/ax
19zIJ4DY6NZsR3NFgkL0gGgp2xQG6imw8+n/IuzRhXATVJtpKvK5iuNwVtbDAhBl5coktG2C4bzQ
dLAMVcpHhRlWPUUBNEBJ1VFjp+5zTPExBmPvqin5epaiJySmLNkD5ydxP+ntXtxNAHbG3K/O/Rgx
9F5KwEa6U2uxuYhyN+9fIOVu6+JFtbgyMmwaoJZRuIGH/ahhZ+NUr1rzSaU4l0Cta46hwsozNrjW
pmBt6rGuPBnh+wYO38LN2Rf7wYsisi+stRSF4G9yH92EeiMZJzOEZd2Y4dtR2bA/+Z0yuVH45T9V
Eg7My1584JVaM89dYwW4AWeywodfC1EcDsuKC+woQEoEmb1wtSyTUJR33CpC3QyW3Ttszza4U2OA
h0UI8T/FCu3TS9f7lMTOJRzt+Xd5uqpNYJdVAELXkaueHSQUymFGHY3HOvI+EaOUCWIu9248VEc9
qIidEuISAS1zpZDv2kBT+3QFZ+qCEiRIfGKazf5sd0RSTM/Uv0UJ31nMGMITCTfjzl1MHgKSSw1+
tKpHji43j7YHKzAWrzQwbZI713FRbWt8c+MJRJPhpm38R5TnwLAaoZQOxJ/HdJvJ4xWlkBM5jp5k
dcdagrNJSpwh1XgfUddeNfOqg4Wqq0PjreKEPlaka0lr0X8/jXF+NpRTzy0+DY3kVGjPqi5GwE66
UsyliEG7oEUzdlk8mnqVZPUWwuCVQD8EAHpkfLJmvvxrrA4doCF2A9pTGq5ggVZTUaj6OjT747cp
bMJymaLW5qhu1lJzQLjNrjO5Fq34a3kYZf9lC+wvE07g6iqcSjFJumoRNSiczEqcAYo1NShXSmJZ
DVSIeuCfHFkUae2uIjJjMaA2JbhYt3sRZqsTah/6PXVORMHasueTzqpgRsesvv2yBwcr+sElilfO
2cbe1No2Y++annNAInRXFrX0oVH22RXoZCo33fKRMmwzTJ82+eCJVwAw8hCfcUpSc0hoCcy/XDz3
7zKIXKD076AKe/miDjjnmtkhUGK/FCYQOXZNhn3d0lDtdSvyUD3Cc2dNdHd3ydmw3WnCKcWvOVyM
wlv+/hr0hagvx6abtbG1PkwNH66BTkwoM+mm2lqsALk50Otwokg2OVueRuGrwRjuxbzXugur34B/
3V9ai3rjcoOeg0XPSfy7uYxs7aHXhFoqeIcqi3PJZ4YCUvcodDck9uXZaTXkrUA2oqq20psfJBcO
qKHUgnbCKq50VnzGLjYVioEcFEioqYugLj34MFw1LhbLhS9JIT0vOfUfdbyBaN+Vdk3iDh6nARR+
cQ4FwpnzxO1qFMWN6/K8GZBgY63ZVAMxpnoJh1cyxwP3PVxg/9XOCwn017Ch3/jT3bX78gISIj86
Tj2WIgJrmaXoEbWT0QxTSdtq7LjpdnURINyU/zcTln6hsK/oJkRh8EcTkR7blx0/9jSzuR5RfXYe
tvJbEIsnjW0RYXOTfwStmgsJrjhccIa0C3rfXPKqGgxnN0lw9rZ9jF8VXzarQ2hKvjdBr9eju2vJ
3+blQhcskcJHPWUSCj/V6k78ed1PWURtLimPaZuXE3Y496EuuJUSam5r7GFGtrUKiWGw3yZel9eY
MdMg0Q1jqWVgaWNDDYJf846wfObGXPLnXNlUDJ4fGh1m5LeCB5i/IzHaQy2CfjwWmONFrU6ctjg7
CXOxO89h5xUAI8Puqrffn0lk9pMXD82hqFuxyHU7uPqE6MHXsOJMHeUMkHdM3jcbQ9D+LBlEkAhJ
9pgwDaRpSqXlVH9MiyFwubrdnp9bhrp7cpYKhpW1+Z3hbEiJbGr1+yf8OQJNusFd9aBs2BFQdp40
7mt5LhLN08DVVXvxqWGPEFrwwLUJmo5Gev56M6uPSpeoI3x3OxTJYKUAGCdodJ9m5KhfZMpGtWEI
kDSS2aWXr73xcwxPHvn294M92mw/74anQwWSXJNsFif5CPxWVcmrc03HLtiRaSThdXReEtA/YN3U
+3hz+dRfP92TmP3ekK8Aqrx/eUxi/1pHkfoo7jrNUvk26Bdo8T1SmKoVxhAfMrwKvIugpSbc+I4+
OGnToeTcYvV/e8hvHQJihUaE6fn6GJedqqeHYFV8AAG3euEvwextGIofezPYx5Mer2N+5yjuX0cg
ivRhxnQNlMCJcM6kc/pL3rkDW1p7Dv7OSyhgRYAl0RGRZHi/BoNmcYmzZnc5A5vrrKFtERMLlCDY
5EWBvgxjaI2xRmPSFpqDGX39HYp/qCsxJP+BlFgFnkrXFXU5ToRdGkR0SMaJgmPgbaAP0W5N37oU
8GQ8yF0Yf44UiZH1q0q1P/aauDQjBPsJHp6X6OOaq2UU15uncDgcXElcDOorpodLfRHj5KbQJVJW
oOWsIQ0CTO8lvhmT4swGk9zE91fOxd5Yh6Z78Jk312IqjKqZKcfngPxNk4zvhj925b/TXf7ms1DZ
iuxQpWlrnQOnOWcylJvggIF8BwYnwImS4Gl1eaeOG5VFtQTyiR9Y6wyTC32pm9FOz2AyZawJCBYc
+6m0/u2fFRb72gePFdndE1qGV4nRnGBTlnEt0tto35oy6RH8q4fuSwkDY+MDXfTsd9mUXvCJ60yk
onA1pGkK7zlgXgb1YKKiMoJlVHzfAgI0UQ58v9hR+JjJ9ZgZxx82h3QJFAm2Zb0AQou8fobKgVqX
zj98OFtwmlwdeWhWd945ym+9G54DfR+ESF2ltH9rancdxwqso97H1t41BPL/JHdND7Y3H1cdvMzG
5xzycEtSL64+xlrECE519JB6bo9clveb5Pv4Z3rT6Nl728Xx4d61bMyoqdxWS9EUmyZZ7iUpY4SX
68yVsFkKA/JVqdbbFR58dzYh8jJKKDxxDsgLn8yXhcpaDYcSwF+lIKWXlAgYBuu4KX/3SqUf9wKf
ITibruHNQNys1+Agh+nYNi3M3cVlDgQQn0yoscqbMyWAk56oukv8dklV9rzCcjukbQYdrxEOKP6L
AWU6VBjgAlzQDXOYbbSvcqvtKW1p0Z9D3ZsWMY8nvro5pw/ROMFdp0uAYvEBdS6S3sZUp082w8DN
rQ3sk4aYxcQ4QEfwDY6xbe9RZ0d8S068SvGXGAq78zMFeOKrISMhYP1U2BdQtd5O1cGN8qO9qMB1
loGlDLzfO0cJLBKLi1NPkoYy1pttujn6ltl+CM/SwVWSYUTFzWn2wf/V2BV3J1mm2XpsrIhUfFdG
ZYKjAYSzRAAj89gv0G3FZULd/L1lw6vcjldJHYDGb9ylLgOAl4wYW32usy7bTyU0nb/Ypab6+vZ7
PJ42Yrdk0mq+ZALpSOp3/m2GMjOtti5Z36IkYWpv+nJ2gZ296+ikrZXyr1SPCHp/opHvIX3rTq06
XvrAaPKnUu3tq4+EMwGiE1YshBLJcYO2zKcytBEgfhGyB3VsWu75yB9X4+1PJYzb+NLQ8rnqvlNp
BAOB9I1KVazrZeFZ4zeF2SfgKBV1QhEuvWqUfCIG3acHLr9Ngx/BXM89CDI8iJ2LHVpmqgDzf0Hp
HyU495wFdNiytX36bJkIGNelwam45qcWbeIaHXrI1hrJHJX8wPZbQ1Sk92KmCBchlD9B3hrnImWN
NhbeMMfb5GSQVt7U7jj1xqttRn3snx/JyV5WhzYfFrimGMhD84bQoRMh9yGvXxeK8u3eQtluiM3g
rdw+OLqQPCaxqIj88U9JjVXuYdn6bUBCnAKjNjw2ml3euBKJ2R9EqO6QFERjFrLNpoNg5Lv7DTT+
gvdGGqP2bsP0FC3Xa16AHNuaSegrEEI3j+5Qj3gvh3rVCbIVpVUYJL6DMNjDfqQ6icR4Mlhp48N7
MrH0FZWCQWAx+XpOlJ+ulKMe/tCVSgVsZVC75v+f/aCMNbetbEWCWx6ygTEfFFcV+slyqnlD+Vpk
tujE6T6UNgbHwk4YqBQtO8GCvdQf5HNyyVOWNQpnxHVqgaPNOH2VdgzRMnXhm3GPHMOpiAiTgy3G
XdWyqVDMVvc9ZvQ/RWqef06eJi0JfiGhXjkYUcSlYu7bQOnDJhLQwEZjA+t4qE88cXNGCnmFmLq5
XRozVKQe3II8Sv8EjuflAtcbXgsTSLT70i4lpj5ibC6S2nSi5mDSvkKb+63WHK/Z0D1CS9NgBadA
AAcQoZAnJbcV59hbL9oURMsd7Qdo+m4Fvh23G6blLqdC1e/rOiD+NLErBuatc1TW2e4/mNU4TKqg
hzL1Xtt44kRDolsBJTDV3vfNqg3GXfRdCUts6hrv8xKQqzlYTs0ucCfLLPadQAznaqyRQOdJFq+a
riC54yat7+4Ak91awJPe47UNN54WONQkta7fc0iYdJz+vnC1LVSrQz5SAn04kzGHhX4XKpvECJf9
3i6nlkClsbksijxB0+KBf/LNyQ02YpufyVz7WJpafHGM2vSVvarWIMM5S+4cK+9iy9yfV27yk52d
/GnNxhdaNDvlgXv4wDuF0mXHxwoynoEcLzJjzQzB2bMiYzGEaAanWEPL37xbNwmyXLwuAr3QB8Bf
r0tjujgc6s/A17k1UY6sWCpduCeIE3l3HIpJQzJxxrgz0V4SJG45nHIlQKtl3cnzWXG6lwYkyDh7
Rj8YTTFWmpS2fFpS55W/nzLleyTq5VSBW+xhTi3ZrFG/he7Srw6OhWB5BYF+fbPHkweFau7nTRBo
zRd0LJLCr9VFAC4JLmlEWFDxYR2kNY0ofM/rrxIhedp7TYDAf9QqFt4qWcFbZtMEfikY17dDbanL
OJxrN0fVyfKjhb4oE/E02nBa9FGmjfImYXLkM2EvrPSwX9n3fPyN9Y7C2Jtjd7oNPjOrniOqiGCs
bpIlVGl1DiA97jjFbvImRTwERuqeIcS+m79hxQpUocY4SMEvclkgJQWvbWMOj7Ogf4NBpgcT1azt
IUohbKRyCo2NJpiKCjeMwWCZ1XkyEWzk9723VK4lhWVHjoLBMCgVt732SXMXoqBrVJfY90oIJ4Gj
BSoOfJEbL82W2cA7kTezSD2KOIenuy4+SvdvcYRtd6gsQEfqVuuOI87WU99sqUBVMhSY+KPeYt+q
t/ul+uelX6+Az3gC2cGgymX96cYt+rGbPafo/dmxgPj7WU+WNXwtT4xvv1Mf++Ni8u/q0T01y9g4
l2GU6X9u/tUA1WvqsLC4nQNP83kA78TovaQ0HoMG9RhpRLj5RxoSJo0LRi5SX/2ZyWvkx7r15UZf
h6pcf4u4W879F4hniTxCZbFN9+dGEBQf9OQrlN6hFQISpfJUmHcjwsgk6LUXuhUGCmGW75yr8HGJ
lKlWMFhHbggBYngBo6c52iiR3pJgtFMVPj529/V0mmGjH5g+hLzuW0EZC/LFDffQ7w0sIhIa7Si3
93C/cVSGRVUBAFCMwG/I2SgGwlPDK93WH01sjDQDLZdNddDwY4YHRdhVgTRuXKbgPpeBnBAzLfIe
QGAFtAfvijhgwFNFQj9dGLNbICNEDyWRa1Ssva64PScqarLNPGtJdnHbad4quoBr/+O9x9rMsLx8
CtZ6JrKAHlc95Lg+NHkI0RRaIfyZ2k9g6xXJ5CMXZTTsq+uVafLFH1O9SpifXksooqFMGwKjVonR
lkWQR7V6Pgfh024aHM1iJNOWLYcnKsnjs9DZxjAX4EhGH28jFZft0HvmzApbYmsLUQ1sJyqsrBcA
poJaMl5D/uIVs59GWdo6bLG3oPWCscDEZtQq/BKJtuh0bo37i8MYbhZxhnXfYD3VAfz9Uj9T3zsP
hGO33L6gnFUkZNVVmW4H8jCttVw5WS9e/DIyuiHmu2rvFFfT5MWtcaJkqQ07ECFxGnd65+NWf+Dt
+cYD0xzzt0u7TfbzFdbnSOLnMlRFZKCBVheSOv+zqKsmrRs0FXgZxLy9BkCYvJuIPvQx/tggzcyG
iblGzQrTflDdvrbTGQI7Gkf/7J5IbabXn8Embl76GRtuLBiSuw2vY7zB0VWSA3szmg4cSqn7phmB
QGVbUTrZ4ZYBHiaeCA5BuiBZ5qomUerdyBg5cG3apFpuyavOF3+8fkaIALGFBkHboR35yRNh2yEZ
yfZQBGsT4o45/DpCuXBg5LH4xQKvFAOXvWmArJwkRIwos5xM3U9cv9eOHEgg8YT7noibCUBWfhU7
p5lcq2U+b6VxgzbNllfvWAEEAQ///U3s5XmQhapiJVa3wCsYPuyzOqtoEEPoceO2gVOh356chIh/
H9VTu7plsPZTAm+xQaVESU/N+7AM2JXhLciXNI+3Giko6sHzdnfgU/Ds2wEhBbC8kYAR3kZD2VYB
lKW9SzJMAo/1814XC32CkeEDvOU7VTnAyBz6pjQoG8HoSaUTFNSvkC3i6u+k6jVDIHOwfqCz0330
Trt+bH2Sf1X1WQ5vJqq0jIqrxem7E+vm+ia/70zIhav0mZrKo2X5Ui5kMGiTMOOiG7VJpPNjtmTl
zwpRcLGsAWdKkUJrHTQgxyQy16XRYLeUNnIK9x2Y8nzeG4Bu4sZWRXohSy55MJ3kT/pU+QJ6ZaSP
dEV6peLfZq2//NACpKyU1HwcRwGRtsTaqQikhjlcXytlKNMiifLOA+Fuyyr6Qis1q7/4yLzlvQ0r
BT+0LBUix3buOx2lkJJoIYUD3UUNBby97kEgnMIqB8EPNSK4F1EmuLmbpMA73ycZUkjMisR0mZPR
k/IX8yM5pZCdwrodMvgw/HKOmh7WofsseEn6W6ogBssfsI0rxZhqvRXS2eoTtr78JcwdBGYesW3L
41tf+BGuFBW6opzNpOcXqdwhDMcH/xS6z9gdEn5RFIiknywjwksER1hZTatVq74JhLpj3f+O79DT
FdhHC8ZVgSJFxe2y4pAJ/XzgUncLtZyyXAySgmIgdQ7cvvUtZDGnJIWjfh8sxpsOv8t1MudDqg9y
D8t+k7ko50+ye/JfMTWV77YdLQcBdCzNJM8lJj6YmjV1JDPbNMF+Cinz9nDiAsrKYsjlI/EOb70Y
r8NA5yz8vLJMeUySn7LlHwfPLAHTT6+4nutoNSO+GNpeSg2Wxfn/VoEZ620PBrI3hvNIzTBRX2Ho
H263vrKsUYe/CptcYuf6T9Q8dZYdwkuY2rcZTfiUoiGWuoNJEhlZX+7DVxbNK2EznqgLc5RjSLrf
hoqGCQNwaJbZuX57voHLeJ/xpfzQ5F+2BgNFkqqweM4Y+BPAc7eqJ+tivuTbZmppFK3QMOOr6LmN
PtlN4LrDQ4dhDJP98KqVBdqPab5EGNlWsAxKAJRBcaGNacEUl0qN2ZK6/Lizr2VSd2E4YfHZ54iD
OsJV/j0VxqaFxOzdj0qVLhEaaoRjQibvMWaY4xmtYyqbd2/45qFPuTm/2M2c4wVyEE51sTXnNFUY
4vHABBXISwawcHruhwX/0AEKsDz4BdGPrxfQlhUdbKg1IfAwZJsuLH6UF8tgHTn3vrEfN02O+tC0
xwaHzpMLEXQtGWN/tmlbwb4raQHF3ggEEnhLp5h1W68dsEu8uLoF+SCZVkfZXIn7aBeYqsuLBagr
354O/e0MF13p2m3vuOfKehvnd4TdwwBrL3t8U2kqpzGGAIwy5Iti3Axf80oCp+b2NKlup6cpMLhH
gye9yaMrNVQVx5HbXVrgbcyfyWX7YJ+RVOGgZoyJoTYofXXslUbY7iWz4KdQI/NitnoFapF8R2K1
NwoFMXSxE5bIKSQlMfOJAWTmSoa1OBMWQI2a7wwK65eFMXDfjBxfhSp/mOe7KWYX9LfGLmF9MlQb
AKd5u/S+pkjoSm7rU+0yvzFDKwmuGPjQON+YNhOUFtvXHP5xuL5tMf+BZ1cmh1kWmUxDKAVZpJmJ
aeYKB2XvGhLAhzv2btWf4+TxaWuxW+jeZShQf0Ju+mwAD4hlIWTDXKVH0K23yITrbfh6Nwgv+FSL
a3ryhHNJviQla8qEsr5/MtNyghHoddwJjNs2OptO8HqCFXaxvXqfIZ2JpbeQ/XZtGWK7hlNsRIgO
JiUlAQVC8FKQr0NHZQZTV1LXD4WGuJJ9N0MNmJQ7siDbFwmBGNBeab3suoPcyVZMv0dvmumfjz+K
n8/cwOFB/jh4D9GHSU51tEoDYjMUdrPVlV1EfcWjmARKPDPFgPM8uzrkuBwQ3dmh2Ymiw+n4Vol2
iBuDGWgKNITBKfKwAutxbdya80uK5/hcSeiQwDwqtFnCniV0mLHqaOyhkYq2MGeX9NspgZdRie/h
FzT2vreKqg2benKwdPwrLNAFvplt3hs/GCtnUczmQ/Hw9O3aB3MYb4ab2LXd1l8u2TbrKY9IWvYB
igT3th2buRdVoDy5iiFAIZ5Z3vlpQmLrhnEwyBcF2V0MJxSTrzQ1Pr9adSISloF4ebbfAZ4QTeXo
6Js+36rvpQ9ULGQsFeeFtFS2Cxiu/ESvjE/DvE5ON4qu5yCVJmmlrE5mI55x9tzPXO9cItd92ykn
bYjAirfyPDHA0YfGQZarvADASE10Nm4l2HbRe2Z/jya++cEkUk3t6zy7gqHeOgr0V2LVdqN7GjkZ
ay7to03ZpNA91scWXodq4iSieAgPtevFkVkU3b22PIfTFdcTaxfbFFzti3oX1terl12u2B6oCawR
kZlXd0Qx0PMYwo3aV7cYkJnmhdVPrC2iyq+3Gi+P+dVfEcEuM4gQsUvqrgV9D7L//w2YoU3fSHmQ
cz3sCdV58l1ocesebVRHh4TL8GgJKjcTb3cml5x0GK3JpMag/0lT82EGj2mqj5h3gb0Tn791hTcW
kY7TTvoqyGfrTl7ndTpjItNPw/t6vDdZ9xJmMNlcLbEOuUt9CICLkqW5t7SJJoKw7zVv3OnrRL/z
q6xK6s/0Oye+0GdDqyyOgHvWMpeZ2inoxjgtR7+BVmpr5gljDp/JMMkTOq4F0kriZzWo/9Hd6eNL
VcSit0qU4tTWsphRSCusXveaQJTIkkeMTKsSjTxvRIR4ZlrUlj83e5W3YC79i32TCcUppqaKrcy9
S90iYkEksBHUINM76hbSDy/5Y6NwqAMzyzG31C7xQXZ5GMpnZuX0nR/iaVP7hZ62KfC9ezEZ4IWf
s+x1NeA1whBsJjfRc3widp8VjUfwxgTzRpeffjr3VQ3MWQF8CDs9vXnV2IzFWC5z9twPKa4YncPo
arfI8RPfqM/a9SL7SzMkGEB1lmHM19CWXw6cU0KjwkiMGbEp7zH8wrtPDvNTVNvYYcgWyIEJxVkd
p5rkXlhNe8PZu6qlpzYGZlEnkO4t72x/d2N7YT3BlHSfdugNjzzz2FkbkhXd0q5F3wlFvYdPzjDr
Ckq5wX2Dx+OAA8hn4z39UwP6ACT70zMLXZaU7h08Oi5Lj3aKYbE5bfaqVuoefTMNQdPvEUI/GBMG
M/ssOEua450FGwcAmWR0CL4Ze58VEvBI/k921OKz4CsulF1sN9Ie9Y02IQ0SLPn8bshbq6Omxrx0
jV6Bsui1oiBpo6OeI63HgIBjmTvlCZxtJ7QYLzfn1UT7tGR8YXLft9IIzpN7MxTBveF9JDbqmEWd
OgEWoZxyoxxqrpVBHUX1ZjLeImaefUDgPEQOW6Veo2dmXI+zVPY55v2n5eyQQMiVXeSKiHuGKCR9
JlANfe+4CPsCg/OGpHkxsQjtgveJvO5gJuve7cnx+ecC1Bt4iEuv2dbrwsZcj8g62HeOzmHY6pyg
Zq70hsyC8zlwnAMJ6xsmeYrfwtxQDBm27UQ9J6ggJCgD8CxRdd9EZ1yuTm6AmmRfx4wv9hU+PPwF
42/vAZpuY9swAHzMkPuD0yAXSbJ/B6TND7jUUJY5cqEv1xv5812PsPngJ71aTTOZZ0hXH2wmsqUy
qTq+VAEW3rLR3iGmggUHwm5TwgeXlyjswpaBjh6g3mi04D5Yq1a0Y4Sc/AePWcPvbfRdJSkVMfsA
FWMp5W+j7ce73HEhaRCS82htiNFCuKcMqqWc7rsV1Eqh1Zgs/yBQanghqV41cnuUWZgVn4NlLhD4
JTGl5XZYqzZ6EMJ5g/+goK8XCL9gJ2SHSCYvIDF3WQjYYtvwpjQkTpT5VvadQy8pbGR9IG8ZgAAf
T1Z65HTxyWkca9L/lMVSlevJafR5WCabuxSLvKPpp/HRlAtJmgX51e+5MHMf1LOzgvyixfQ9o0Tt
3aYOOTbHyHREDrqgP0hb08XCdorYvOi0l1LK6N7ICKtxgC+nEYXZY1hzXmRUHzXlRyIyFcYiZRui
wbYpis+oPTQ1Zxm2soHH0hq91B78gaH4tlh/yOh9CV9NQ+l2EyivhyXkEmiisn0lDZ5DOT4W/uY6
HNx1pMELGYC0Ohbr5TX8K+XNUpXtUTcCglyzbc/ei6FQnMNkAqf0+gzwQ7hX2uIR+MMyp1nmC/iw
t9FZk7P4SKpBT3IdjFfcqEUc/QYx4yYQwzLPspbBqVcXaHeVh6FqMS0PyWNatR8OjQXMC2TMSqZ9
2FsrNUV+O47k6PEAinTTq35NcdnTRZO3R2vBpdOSgQs5Wkjt0oxRmUF7wLzqRoPWbzwR44184Qcz
q17H4BkEnutsRoBGero1x9OyetpREZODUrUtFdA1O0nYoBqgI9xoMo0Pb3TxmvOSi7T14LiR61om
wU/CK41qZxW80IaPUr1n3eS7a3x8xDn7khnFKCjKPsYxm9bxgLOYI83RNMsJ7i6tmD3+5D4KRmSa
8nTAzjAZEKs9z08Es0xboPnze2+iDtEhF1hhUiP7kHtByIMg0JMuUL3uZfBnKI8Gq4ZHI/MeK9//
qgV7vr7XxvBHoVhOjVcAby4Aa9YKRqD4KYiC5KpQIG2JO46riihW1e98k5Gg0+XYFXwyyrpxKXUJ
uYsV7IMnULuRLzCnJYhSW82kUa1wBkeiOsxLb0KCMJMrCvnWxHuuNUdwbn9SdMw+GckGVPDkaj3k
8X6zc4HK42biDR2fWL06C1QrVxqbcsD2+T1Rbq72hQdqvS08Qh4Pu7pKQHuzqX9NZaMvyMtvFco0
vS+LzgKkAZUAEbmF7Wgpr8r7cZWATX6MEyAZomaEDWM5EdnF6t8CnsjMmuM+3e+tprAPEtfkU6xZ
gVd8dcS+OSw/tdoEoIaERMZ+TwA4bl5DAnmdtwGGiHJ7KjBYacrintYKO1WGhv0cBu6J83JzWqWK
jsQZbGBtswOkyClVdISXLKCfGwgdZqBVSooKfE3T+oDHXHrQU4FfgUGfR4+jAir+zjg9mvpsB65t
aWiZHH9AdF5j6QSNGZzii4/qqtyRjkHK46VkT2/9cpD368WShC6haZqiAT/BJxqw7Qi/MJ9zenue
SufBQXXmJ7Ybt1clyQcSxODgaIXHUwHjHAtQA3pn/XmK7pdRluAMj2JI+MrH7VyJls7xhEbznwwx
rxIKHDWy5zhAhNGsMSngO5x2N6tzvz77MYHjiUHi+rB5CV+KPFENSSzjrDX1DcqKGxO9UFvzdQxV
qJBK1eqeBgFyf2TY3F6HIDU/ClCqU5I6zTBLfxDZPoFh0synBxrXpx5ICFAHYEHMF7r2MZQa1hqK
53KRzL+RmWX808ICqXfA7Y2rXwWY7tbNN7tmGju5A4aN/ny7mj+qZd0ERif/Radi71cWLUBKBL4d
dgdvdEjWenPTeKmtAIMsqJabTIYJSPV4q4IOkUNnmJrLUQXenSmku9r+O7wdJBSs+CyIeacdPiHP
rgCQDvDQ8ZFvF4vZYRx6u4rQM1OhaWxrnWCX94bZiYuE5Bh3mHU4gaXS6fM+rbWPhwVUpxILEJJd
pUYR5Y+7XXbAv/FeDGjvzcks+fF9Ko1huLRf3Jai7qz/D8nMjB80TZGIfHiZQJeMpQ/YO5fvm881
NVHjJBFg+z9R9xsVORWgahbO+09mDU8h4liN8UTQIcjNR9Iy1laTwTQuHzjDPQmRUTiuGVoQc2rW
omxOQctfLc9O5StLt2BzOyDeQ7G8j2rT19hBluIzyaMCnfbAH8a/YHOQahh90eQcKLmKwcWocw1v
yCsq3/bpIVsAeAfv6ljT1t8a8kNoHgnCueK7AFPtU53WnbwBu0NomjfX8Bu3jCUwYZCSja5kMHf5
Rh/B01h517j8dsAQgOstMtdoI74FmSPL0yhrcjzo/NvH5VEBo9pws49U8ZH0fPVCDE/3BoWadh3M
SUosgGyf1IWoVCx6HzCXN4qs4ucaTMy/N3FUuY/lDtGFbPudDxEc0cbn52BBnp0rQanYtgYHp1K5
CNUIoHUSUwlirrfoDbAUalJh+o3rfFEi51fbXPWjIz0HAH8ibDq/0fBn4fHX1eDroU7jGwriTOq9
GOSwdpAtBs3x1905Z+j6Woln/uL6oE9SVwSo22+L3zbGNJg8OSma551L9N4G70g/vPYUb5QbJTpv
TWnEtUXkd1OdAnx8b5zPrVHaxWbCBJpMbHQL2TiTzf7Mdf9IP2K2FpsIpHm3xJ0sUHtylFFQF9Oa
3Ors/WMubPU1qQ8vRVv+LfuYleLBIeySnDZisT5NjTK8BCqrWlO7Hqv9lCF3R2f0xofuUEMargVL
b0VG96dwFSCL2g/KxiZ3kOeOh6xy/IPJiruYY3KSEeFddvMwLwP9mVIujT1Xlpkne2Imfdmo2Z8T
azNWsqwY0WrIaZ5ltsGFOOJNmmMlruc3Pv0Li3zraOo/VzHTmgn7Hd1jE+tVawm71aNB+zD67qjK
wEVdJNgB0Q3QS8h3Jpd6z6tTsLk2TyCBpO8saRZ0wSXppBeOXpK2/7L9dNkca7OUULSM3BUvoFvK
po5s2WiX9SlNZEoTKh20/QRwWj+aVWVhJW0w4QXPGcveDUkrXbGR7mY3OOF/o11dqdf0nGuUpW2O
saXO0jtgZOpC4pYy1NfGxL463u6gn6Zc1Q9a9H9tUcMY5NW9NZTa9a/ziz3ThJC5HIYktZJTCtgX
FcKSMJYnqZyKziZF5Stoej48j3j/vPm7/7DPZMYTiQlZpVFhNhZgjrEF+UqXPlDfYkdNTHnaK770
W4Q4hSrEEijlaZeN5lfyqjqKPAvVnCPlpJ1FQGGWTJq3qzQBQskem92XHJmrgDQidY0EzYOKnyHn
GuBffbkYj6YaKEeGWQJwI0IWuyIyHWdL3ferP7TNogFSRk/CkKhjRsI9Hn4O+b3AaA88teZW8NAF
LiNRkNsY98w2onmMRGqFkYG1Eud8X2FWWnxwP2+BPIWUYgB5HDYT2sAxDeDGGJXF+rTyppvGYoEc
Jn11xM/quy3DWCVaZs52Y6fgerzIsDJdHYoX+KoNjIX4md0POzdR6JQPvHBM2G9lFJGq3wt+8G/A
KuF18IGBOXW7Y5Hft1aT225kL+y291N+0tBRphym9cdhCejnXEUF7PeYNxY37FwqGhVwZc373ynw
AND+O3c3+AszWfL/Jwv55CLUidRhktR+6PQh0nA57pq1et8VCy06qry4WISzN5pxcV7bRtl/vAPC
Vrv6La0dceYErbsOEOBbUymMrXySOb1hqWJ/W4kIXXgZhn5xASSLIxTUUmfAdHU25LHCy5ikymD/
WAt+7MtUk6G1GmA9UASSDReHl52laFI2opD1at3RDNbwZhiVTGhq864LB9hPtmUYqYjEeY3b/Evk
hT9RHdmQ4EwBUD84ro6STbEsMShn8rOIsHF724gdf3CoGqMUC6QHmDJUiXj478ZPmfLpkMSHW9oh
WH2ZR1pg6y18QDz/Au0FehLL7qmzuXjQnepSsHUd84KOX7ftdCZmFcPl9msw077czLhjrbRmE3ZE
QnjAhuI0WJXlMhNuVf4Y8dpHv9sOKUyV/1U+Z3HJrfl711TPCTTeUP/9c0WAuMoZlyU43RwiLLhJ
2kkoCyvcfJgsaKsURtK9WGSu631jHdlTnx0kNis3BMn5ZoD2yvo91ysmYRj6eG2/9GyOGkWPctlt
NOolSVWtOykN4hO0I8+Pin6y0jnKZd0Byvy4CXJD69aD8Tf9pCjwBsM+SiDMtem/9srDD6tyhVXU
272y2RN/Of58vJ5UI2TR7DocPh3QpWSQbBVcAqNjEw588MlJ1mAAh/rTNStSmPNpTWjkRrywWKFW
cyNW/i2WYK3KnEZ+HAFC7ouYyYRoicMk1JvFlwRVmFCNOzStWpB5NnMU9eVT4/R1ZfdyeyPAcW3W
QAbIVkq2s7YM0tfhHSBBiCFynNcZVHSJNrneMax8RuBoZC6OSqxGDMo/8UF5aU2uIJO0+egaX8Sa
okkXlEBeLf+0yz5PCkzQnJf9Ahvhgz7uRnWmJ7KhY+2/c6exHqs7rXVeDpvxNRP6fvXb57vORA8o
KHC5FTscRkScKHdnVe9fdl3Wd7AsK7GSaoe7GZ0/o/LtlApEfjQhbQturGJLeQXxb5FtaLlHtZQh
wpJRPAf98xsazjh9ICcvecFl7sdRLW5PRS8TlD25bC3zGe9LrpvoEUcqtUoX4X9D8DtEzvsaGOPx
A6N29MLUByl7ALTz7Lj7eYrlRmSDr01LL21l29r25hGHZNUoIcCY9aXQrq+tioRqFBkY0a6mevxX
bKEdgWRV/OHUN1DtkQszSb4HQN/J9qOvA5BlAm72SeNtSXpIs1X/l2ex/69kLqdocOgqHhKI5y+N
Q/uYqmpAiCktNKrr8F+MHIrsFaqxitjyCvKGuixDk3YNsGX39vmCJMPdtJgjYIasZ2HudGIU4HBe
fV+o6Hsk4uAz5CJgeL4tDvwQqHCct1CtbcsnFVjb0071dDMwqKHRSCaTCU61rJAkRBPIoAXpKl3L
znxKyX9sRfKFxD6wgk5xR1EY6xEbdw+Ld4yj54ANbspuJYZ3qYqEoVSV/CjP2Xj9hCmvVwj6rseZ
XVSUfXiGjiX3AciSCuyjxleauWuS3BHSwsdRU+RaJNH2kby590oTlg9saK0yFR1UeKhwK1jt74JP
piNsuofa/Wmmlbp7/CfpOQ+aDsK+hWDh7qIFx2FqSP2S/XBsVDqlCREcnFBhGTimzgayJoV5A0Gv
2zjfTydnt9VrfYOEfHg/raOaxERbrEz95Gywu2QICn9TqTaRB32M7tmyx141SBJ/Z05W8Y9lYlYb
rx7GnUiPFUIx6YGoyXF/oZRV0kKfL2f1Ydbgf086dbbxjPjVUT72+tOopNPm3pQ41JhgjkPdn8yF
aKYsgwF9GJfbEIRCOdfSA7nP+Soyz2CRwqIm83BRqHwbi2+Iy4IWXWhQdvsfX//Ek82SdrvMua73
zT4IOTNtmr/FPfOFwobU9d306jX9qINbk/7OKWf40w7pPB8sIU8nV0CAaaYOC5KANviDrZv5azeY
XGwxHFWE1yF43BNrCcGvSDB0u3bukW7ZMD0ValSXVnaCs3wZRq7/QH9W9CxfDCDnhnZYF8wz+EYC
Kb03P8x03Rjl/uqqyy/XiaqmEs/d81J0Mr3oe+/q3KQhNbQ47Z38GPhJe+AYqzr5rtHSo0g5H0Yi
uwjc1hWltZMdiNexvb1hyXv8nCZIwI+jsHPqGoXu/brLPcmiUF22dbGita/6bvNbZ95tyvOY19S8
n4h3K7i6EdGrrgLF5VgUF0j8IDRU8UDfqIjmMKfWWBpgN4joaWsxQqo6Nh3nrxKVbTynoMuF18lB
RLPxHLBleCvtwfUtdrrJa/bhBOE/nIykQ4ddP+2VbdtjrUWwL81xYfi81MtotWoLhENXPKnVVszg
yslIZT7kL6j+CA2ahJbfmJRw5yHchpXaEREjXhPnGW7qIRaUUjPM/8G6WlCNMqXNY40WhnsEGK9n
6bUxlvHUgsFxd7l8BLPagiVvmLcuD2l9o6nREexV613U2KEiaqQEVmqFdzHeH2aH1gxHKd/DWXUy
r0872Xa3kyy3H/gni75wCD9ATsZMfuL+ihNptCz7iE0To/Um3Acg5+C4HRMVYeDoF+4f8N8RQwEe
RV6BaSX/PwI1J3Yr/QxXhGiXrcHhyhm9jlJ1m4COAvZmiQ0AlvLjz1pqe9naXll7A5uOa7Zr8VXs
lnZT/U7Aq8z+2b539x6iUHocepfzo9uX7/L8AmkHowL8XaP88WMk0Wk5a/B2w832ulD/eNlWNATn
q94WHR0BX2TrNtWCgdMNvpOTFulkpDV43AdBohyH7mGSjUMLiUMw9mzWfjVQ5HfB+u0c1fbd1MwM
u9/XohgbxyMSzoRRFtJSTtG2Il3FFGnjHm6tyw4Z8QmTaXBI1ev4xf0IBuYsl+H7PqzmdhSPQ9zG
KmSNNysDbmlcHfhCN9EFJ11HGB1cBLg4aDa5Xv4M11xjTSFoB18Ta6+chFxOdkz/AgjV5iH4D2HA
G6egaYZpvMbeq0c64QCSS1lRi+FAr9QIV5DDaYNSFQXvYhGFkZMrFp1KygeT9Y/4qpisqwOVq7hn
uwIQKM7z8QQULRJcNHP7EIJhcebgCoJHgrH3wIzKgXMl931AmDXrUUFJeQWJYqa/RkXazVcZGnYK
p01a1eWFn8fblOwm/EJXFpcR2A8SE0OqmYwji/KYb/dmRHpaWrtMZipflEFObIQGo27NghKiS47o
rbnph5/5lI7+1DiVvaBPQMVnt6RMaqOlJ/ALIQu6OkSJSSNB7nikimxrTs7WDW6sFRTS2JlADtQA
FcZ36BvNWzAwmTwfoaMxbw4N7uerfkruIn6QKu5Io83LwKI26i1kh4Qgi5HrplR1ylpd/y2hM47m
elt5Jwg+R9Rj0gzfGx1xyfGVf5DDQqfgAxzdb2URd8tTqt6REoASVKTbJYFVSz8lFv79iMv+dK/o
DVlvfQQwFzOuYAzoYqHsOskTnaP4NvPoWXM3+YcYuBf94Tp/wE2Zrwge6+ZZZKpNTK80yKkW4fqq
FyW1vL+kfhHWV3zmjchotdAiRNpGu9Nx9a5c0JBafkrjNed7vBwZ6BWK1JbBpTIF0ZJwy/X0ikEt
VGfNJIPTWJyXQvBxZyzkof6v0W5kPZUbn+rau1a0k3voN6HVvAVeksqo5h/BASGwjS7RAG6l3ENP
t/LBvBb3xIILiE/6G7l1U8o0k0PJY5wiHdBjER1S3j1+bDb1456wcJEtWrr0qjcqD5Lc4uBVI6FG
GhFqeD2fwT36tGW2NdHsYJBLbuWI2atTAa5PdlZwewoZ/dRCndCd3LyPMV+8X/Y3ssub965NFhCp
ktZQJdPR5rOGWrAyRpKroelRASFPTpOlxa+e3nHaVZ9eOovkT9WxvifbPizxnlk/bRUiYGiv0R6s
eOk5gI62PmEbuGm6oepph9DhYiKqDkUGPsesdhYCPM/SFLIQ7xk649srXJ7V+6/I8IrVQVy/pKZh
b+zb3M5sHjfWK5CGcFpMdWfeQDUzDwzoCpsD+9DDTFgUUhGCL+zl/Kue6RP4pPHFdV6/zy+F8fWD
F18/S25WBpy+pCQYyLkDsb5M7n1gi7lQnYQ3YY+HXJnQjYdt+amspPZx2ke1azYE7mJ7EWeYj64X
nUz3xKVm64TB0hOsisjcjf49W1K6r3h3JuMvdraTFwEtUqqHbp8ix4T/gfcngyuyWvBiOxKRXbBt
TpblPpCwq6i9QQf9hcvPLo3Yc/XU3Ug1+0xKEmZLmqtCfA3le8/NSraaQxU8zvKtvflTenvFU8x/
T0cKdbxPzDKJkS6MJNx183fuXHx1X0RDgAiSGLceLS7vgoYJofQSQs/zEU3FoRAu+pJ4OHXKkKC7
aYxpzYogeFflbSWw5vgOGzrjdeAYbRtj2EUNFusXLPDyUzBWfIeozomIaTFpOjIlDUe8DfLtehsL
iTjd4lcnsRNBkUTBbbO1/p3C1+kxhKTt7o+WSQDvoYbeswWJnz4lJw9lLYrv0T7c4r8eyN+OVZCT
LDHENPV3/+ienzgNN27ZhuUqSpyutajBZaDy/5pIFJ7I+SKbutDHaJUDLdaXflK7E0WPnNgilyiC
VKbrRvEIjxSFg3SUWFaJhddh1H+Lr/jIbs8wUAb5rcESVcXEyeMlbBEjVWYu23V69xTsKnkPqzDl
P8NoAU1fIdda51xOCVZqckYs4Gs2w5aECYTWeg11UhTOQ+Z4AMlxpD69g4n3Acn1bAz9ZAfOVl6o
SgG6SXbI7YKORgSy+pATWXFv+LbnbS2DQEB2YCifeEERSGOVgoAfa4R8kwH2kEfWXZwj81CqRI21
hpIX5w3Re1DbNik+LjeW8noK+V8SXO0rVuan7yO3qEhHtOlTBQ6gtd1PLrSG2Guay2Rzxh8LRZi6
4nZduIWQOlk3803xpKk108aqzJtv6+nghPfU6I6EsIsBVnDn/FO5DDa2D79gkUZEx46RBXt8DfsK
l9/9LJHq240azcAEboVY4DzmTlvZkjM3uw8DBqXtuHbu2tfp5mTbatSpJfnne9/W2ZfQaIsD58/v
q9ziGvhlcxUKVZL3r0pLkXONZ3TX6hJJrj7Y4eLlrKWFCCN1LrzhisesckBqJA1NHgPv8xxTgqBJ
YzCtL9k0SMiank3vzBEmaPx1bWbHoeg8IDNPq3M1C27vhsx0iRZZwONbZsrAJUqUqXPHc76vOLap
QrLdsRrHFoCH8RJ7qe12yHGR63Q9rJYglbDr6scuk0YYoJDqP+ctTe373x8kU0DvhUBnh0dFbiBI
huFniVdu3zCI3KIKO3EQXiN398j3o9LXJE9QXUKFW/uRAvg/IBmyHkdWJkWDkcEpPgzspKEfMN0B
PKa1DeTgj3rYj7X8JTTzCauLdrlY+c+mtxDnAND3j8gySH6mXjXJnJM6jVoX8RXk8ZFthP1UjLlu
nFvFWbijXbyBc7kyzTXGOhN1xyPbu1bxQaEQWe4wdoqMI4wcRn/fO+gJ9EPgvJeON3q6rYkUWn7V
iALniPy7nDrjw9DEi6iP0beh8D9NAxdvz+TKGmj4LXvYJ9krLOYVJPTmCCIrRCfUxT2+WIGi6AhJ
+mdfwbOYEoR0zJmOMR9+NdduToFFxOlBOCtoqCpEztC0+msarE8h9B6Mmj0IolQpMdx19glJ3BNj
I9xNgSpvg4CyQjjaDQp4Ql/jQB1F8Xl04su6dkIlnl4PV7SzV5Cu/Zu8D2Oq1iHR6GtkQSA1m4tO
jUrN7D6Jx3h0nNKBT4ip2BmCU+RAO2FfjSHl1kDcfEhyX4vMiWvl7XN/ilNEJadcdg/CuscyOyT8
iBa46NFC0L3DPxx9CjF66tELJFEokxhG9MhyjC/MbYCN9sEyiOHXMgEj18/RVbBRwHftTL8zIgsV
K4AxcLicowTRzroNU3SNgrFvt+EZygmE8v/utSisD6tW6mzWnddGQnjzsDU8IpjIlzuoOvU2upfP
YDtOxJW62A1/gCqTZoz37d4cQHvxiXJFxcDIwZigi1o3HjdM9aG4627JO0nbvUezn6w3bjXCzTdW
z5mSXsVtpnsD0IN6XtHSl9Zj39OdZnfSGRy7LU32lPdHzRJMyjjpC0hudT/mcoNuYXEvxQ5dw9yc
fgsHgPlQAUcJ3GFQ03conTzwIx9bZcIxmR49P7wUNZxeQIKoalbvWvsUOrMh+46zoTdViqok/+dy
JKoReKRG+1q6S2cFPmKOdKpBkuSAjmJ8J1kdZCJF43bhRfx4LNJTEAMIn0PxgrWyIQI9vp7IS1ud
u4vPDzF6u+583V5EOFr5n2Hz6GDB/Ls/iIMHceR0lhq0frjAmaZzKvTpp4pX6HflglGPR+x2dJZF
qyo4nxkfcV65FUZA/QgfUsj/Q8TeK3AJiy1uTmSyYWZS9tRAOneZqU5dIeKz8kCG88NK8yYRjIcp
8BNlNtjs08E/Yki7ur6DrDDx3mbR+ofL/5CANxcDxD3OWAMLj0kL/oUhYYgBY55VutvK5Zg+03Z0
nr0l6Y/ta4XvCiDlCugpUSf3xQPMfKDp0YTW3pLEj7R1Z+7XB7nqAbDTW3btqb8ayCZI84nEJCBu
LB59hYFjA7+uV92lCg1CAMnPNfofiYIhyJn8hm7bAfp7dr4uHqRYaSdsuMixCbllElh5bjcunrPh
ACaRU5nyrZtM2WBp6HdNJ9Q/eG+wdEce+aWEns+ojQ8GQID71+xflK6sl9j47yMO+avU9UTyb2X/
VjjIVBlqzv6Q+zHMjUK0offsPmQsqEds9rYrllaS3yiefhzuzaYAZLv2PaAkd1nmWevfP4k6DAZE
D1hfpEoWItl1cI2Feva485EUqNI7mzjYi+IotA1xPhbmI93LfIxJ1PU4xmTicABXb1yUj0tpJj+0
9W2Wywc8+N525gB93PWVg96v/GAY2oXG1cDj4TSaKKaeRLOGRSq73ZCM0VwjRigxH9KeK4pssCVV
o8w3iQNdjQ+SilBEFVBN0DDGN4uljvmK8w5FOLtn1T8zL9Cv8GMr1sdG9Artr3FCKPxVhftLCo17
cVCE7nfHbKpQDIaqczWtFIv9H87JLZXcs2Wejv8YyyTBBmMsXIFSS2a7v+RL+sECHOEw5i5Yo/4H
sXFOLPglt8EBrItwHaYiPvANnGNXAMhHwRphAAo+hrpeEI1b9ZchkK/gZuhw7ZMzJ1/SuzrSTRc6
it+L3TZaUwMghUjU0JuedLNKhp4PYXg9QPCSChsJv+BiDAHPTDwUfI8vsD7Pna4lgHfOZY0N8DHr
DwbOsdV0XtGGdnuQ2XiMcS65KEOodxIv2B9IgBpWNeegOc/A4ISuxraE3Ulro6RIRTGWKLo/gHzx
msQWwARDwgHmbLpSpOH+VxvrNzIoIJPZA709646MYvKYdroEODN9PRtmMKKI81CzJX02znwQxptj
8rX1hzQvN3GgU/6QUxyzhgGiG+SlDhSIjqi0OIGk+bjCfFaZdVLNMGwuoZbnWcnkx6rfGD3u+LFl
GPdfl21iXj1zhRNECwmMlvhRUpoZ9U0R26vXlDF+JzrPjBSGIolJFC+7OVvVuLY+GwdOrFxiX+ZG
uOJiLSjyO6pEoYJct5vswY6MTIEaKtMQh9Vc9DXbDWWNQAl2LQsRu2yBj0wzmdfUoP+pUa95XO6W
T/Gh79+JSCzqQBgESkYTwqw2nP3C54EKBn21PglTRjhCOfhYYuBBzxaKpUInAUOQfH4op4JIZRN7
RTdSPO6+4AiUm6HrkExYQG9+ucyq4drHGkELVa0vLb8Jy/9HbOdmB8p0QQJ9CcwLoQP74okdZVfU
Q9ylP3vD1AbLngWRFR4JHJt1HZ9M+eDj3lr0rX0AJKKKjacmq48pk+lWmXGbbcf/nqp37vp/e7Fa
BPkzoENSB3bC6lBvHTylwI1/GJFzpLEYzkTNcp7DXrp63TzmT1lJovFuAtzu/7bFWA5hzWZ4cGrW
W/GfiiMzhnNRNycA1Jub7+IUMnZx2I6mbSLltqmBk94zv9BzUnuPnpTeuLHO3TT+fIu5yluRdM24
DLvSWuoad6WF6pUrSdGxVwm5zNJNy59NCUmdlfaAPw9ti3gTV7giDUUl5QHNVAzBFzSaTXK6WQjB
etd3Rs8aFWa57zdg3bv4vhA0AMIQ93IBynI6x1nyiWULwRVtNhvbu/0gJ3yQsauIKihjXNcaDFNJ
W+jCI0SGNqPcGPl2x2DUi/Uaek/jkVpVXjrs7oeMu0L/1DOmAmY3iL8MH7c9oJyDzYrGElywU6gf
TfQH2MV5iLYp4yypZAGVuI/aGfM9Y0N7+3Q8/jWBPm+AKg/PGK31ckZPXCIP2siXDkb6ThRaTfih
scC+BFQLD2tejCBrwN8auIxmx818xvQbypBbUSvCfycWVieEVIYRrAKT0wgX5taYyOW2I2yZHUZC
cxYcj+oM0/7Faklby6nInCPhXmS1IjrIWLndVR+wtFyg57HHTh9l3wt2RmEGqKv7k/sQDoipafkc
du6pqXtjr3qFmDskcIclC6F28xsosgiApVjWvaOqDTCdRUpTWxcocjJfohcykDbgso/vR7KSxYm3
pH+LhroI5+rEIPhgra4bQpqDDXU5GnN9fyKUxaeH4Q7mP7fCksSfmY7y5uaZv5ECnk3dUx/Pct85
gJzEnL3clTAOi4WF4p2kRYMo1feszcE3ga/NwZ6PATkzcyqGcaQRV4hJsOxkYItqAjg/+Vzv9QQ/
b0JYvEFkVZ3S2Y+ZPuNl8pHo5pp0lz3snJY7gWMrY/+ANXAb6wbhU+JDHydSzZyi4n7Sm/ZijOzs
wAiNu8ni1NVCZ5aXSFPIzyGgwsyQgT9/uckmQItTCpDsH39noXJ9SdubPeRu7z2YeSeU1bZCtQjJ
BW/vK9y+GlUDpJJfgMjvcDqbS2stNK8p18pxnfNf1JCRs2TlQyHTCnh53QFEjJxaaF0gom1fg888
Itox/6SiIe998Prn1W2CHuHLOhhRbInLhrRWyQHl6iJodryp9LydIUUir9GY2H8kRiccv52a9193
zkW/FSF0hKpeztL7NskZT9ai1tP4kKiRL9vopy7nfHy/OjVoUXOuGhKejlAd+jtStah3i482J4WQ
4CBnAErGFn17CMV+m5V9IM7t+C/R10YuFAZXFEjiSpu9OQ1AdFsq4L/1fCmqWv7OYkr4vLN6E11j
v247G1pQLoGv8V65KTf+Rs0dOUtWjcNDCwC6cAsl4Ppk6LP95DRQF+ZqPTxUYcDl4L9zEi896nYA
herSeBQvlb2bAxOC3pbpeMV19L5o8BS3JnIdNJjG7NNo6PhQKtaHpw8DvEIt/SHX06U/cBlVm8gk
FX34VWPDvXlPU58w5PEp4V90wB1DBfPC+7axXojwlIP2ByMrgZgu0Jif6cQatFc50G67VruawQPv
wUet9qVqYNLpGeQ6ujFSzQ8Zgz8lJTcv5ceGtZ7/2pa5ABR6Rpmy9SuC5wZl33jTldBsS3B7PgbH
FqL4y2Uf2Lf8yRnm2UJN7Gk7OizUtn1Sa9SanegIwXeGKCOrnhfc3AEmuIy56oFifgZHfLV2BTPZ
Z4h7r8Zfrs2hZMYFf9M61KiAn0Rts2Ee5yGEgzO4fTkZo77azfKRyhKjjOPgT0HagczRCoH6xMmJ
IbflAEmZQ14li8Er6DTBgWLn2sCeiR8I+e4kd92GATE89gpHCMq5Z0/Mw3yQCBXwD3FyZ0tSgoVA
L3wEQIsG7Thr2LV5iy0Aqvht+jzMalW118r3ZBx65233EFkJKypoMTr37B06I10lRS4Dn67ZIvGl
hIkRXhaMXTPrg2/QcCGyT4t92JaqQ80CV6iCbcIa5EgY1hGP2iKMytsH4T/0MfYorZU8dUKTJfBR
DnT/83vpE4QLvTR17QjFkKEjiafYWBTH4OQOJYuXRM2ZGkD1qdcuEXoq9Z4o7riJxCT33/OQqxl+
NhtFOSvqpKth335jryoj0T0I6EPAQFjPK12ba0F/7EiQZf2ijopQXxJhzbOKj5Lz+N9knM7CII9C
Xg2Z6m44OkuTX7pZDSwoWwkpw8CP4EYhZt2HxwaZIReBFweb38FDF9JoAJAXywJn9D3fq5ZFBRTU
EaGX9OJVXaaMhhQMb/+iLTrsLWo5GJ4t0SzvXEocU/9FJCyb5UfNneprCVjdNp7uFIaXG0TjXBT3
xIXKRKHM/dIpWG/4Q8V90z+6EnAcCETXBocgk0aLmqiKsNqUFAfL4wBZ2G8UAaQDS+9UFKsS4ow3
uECkZlPHoKF6lVmRDZiKoSVmJVRx1YJCJGzCckqah98uI+fQK/GNhRflUsrL22S2p645q+RGfLSX
hwBj0vFYOPZfp09VNjopGGnFSwRiCjp6I5QsF2Ub3mDPx5jyYfe5i9zVq8D0XEyGPG6EeMIVcOlG
4p0m9LM75mB/n6QjBXQE7qfMZ8ijUbBbeh5QZ3P9Q78JAuYxG9I6xVbFkmwmAIkFGgH82cquacxp
yQX88CWrhQcBP4fitnhR6wfgg+Pqwlvlcg5anYMx5dyhYKon3avfT2avgNFzO7beaoUuIZtVIpuT
q8VMu2ZiPWA+H2pbeDYyQVX9RMsemqkNnHLhh8g+EX4RSfE3ilzrTcUYuMnSyMS8G8q4mnajf2C1
fo9dTQygDGn8354c8OSG8XYEI1/dqFBqFd/+jWaJGkM/EfNqaTjL4O6c+fDk5ttqDBWCPU3uEgFV
VaGZtQmWdYcbGOdxQijsm7456uBN1S+K2Xfl4fmqQgUnIn0azW3ONrTqNlgiHby3aAOVGvUELSbA
vNAXlYmzbGAmFDlqPhQvmsWa/I0n/znLswLGHdylxym8TXZJUpeSkrt1zckZDA+3DlfRN96964sX
yJrNmlcY5pHRfBOz2nHDKj/n+t1hqv4BcwpqJRCJWg2n/2imm+QbeR3LbWCzhspuOT9+NuxGMcfv
a9RPRXWMqhVLG676wfXlbB56iRn3FQ5PikkjkmeP0etLEbAj8ZzWBqN+k2HQMolUOIiZ+SMo+RNg
ynGKJb0l35Hcbhye2wBOIHBsHvsWM8oLuWmYEbyaZ0yUeSMGNdm8LGjPwG1J7q7BXkxDty6F/+Fu
aGmzUwksFdHRLhOXOEOib5wRSe+PHgOsJqk0fBghbrrhZTwkZy9s2rSHi7TF49e8yHxXpRa32px2
lb+MLJEQ6zR5j/Dl5UtIoE9pKQdDBoXBnYZdgowrr/w1q9maptjLzpsa9Fs+UNNSEX8ahZ6qk8/Z
uG07MIvDmsqb9xpbbb9jq1kJTGerG7b7as0rAIVrLNHR/ue7bTwdHyWstvRJZzns9VhmSctt/7OM
SGDHK3iBM1V+f/VrIOGPYK8sSEMR6kMpxk4yzU9mHnAudCVMaVDPphLFMObXZJQxTHYwOKYdK0W+
yPi571a/syY5jrtm2DZWt1G7ctGIHhYmTPxvT3blYY8trizb9LQt7xDdlNc0n/R2A2EtMPkxIrRv
RC7BqRzqcwIRJ8Wizjio8rzMs2t+RiG2iJO+uSRancQkhw0Pc9+pl2gGztAD/aMWWx3RDqb1BS4s
WE0CMOCFrzycjbms1vXs3E2pkq+k8AkK933xNFjdBXLsdzq/CVYnDTe/pHL/UmvJSXgaEMW42eYL
gqZO6lmWn0MoVd4f/9RYQ1Do6/F56Yw7q04W2IykWMGzfg2eTAQbBjdOCn4FO9xQvedsXlftXx8g
DeYga04ir9lYEGfRUukWHVTnwyJ3JgUAY3AWo99hkDRkWMCifTA2NigQQPKpZhXbEqez8cYs5e81
drmcmqI801CCNXfphAxyaVOaw08bfREQDfYd10GrvDNTfCR2iQkwe2nXUkhXkl6sVxVmc32N9FLo
x0bExohqBPTJfZSbMQupm4dhPKcMz/wxLiQYBvLY+4PIpW1vs/VYPUMgOoNHms9h5/IePZfJAuTR
hKq6S7t9UV/Fbj+vw8adXFRiraLcllIHqSwOrsVhH7xrFu4OWuMxfsCTwKEKxAh46pXO/MjPu/Pc
hg7jZbC55tulHiFRiwMQipihnhhLRQyOqcmTwUgbyiCK8fdMvp3eYzZx9wxlkC5zpLQDH1yV+Qh3
nWXWdJBy3e1PH2tRA2YpVWeSBRRAC2STKpyGD15ullHT/NvJi3QXnethmaSz+fTvF7SmALve4Ptv
eF/NyF4H7YksGkYrFvC+hxQ5jDAX9IUE32tbqltKt4D5bWUjZy/NgQIOiDQow/XtkwVQslBWLXeo
IOKYLwlG0weoPRTMof9fHWoCnclLdF9FpJFUVQP1Z/gWdj8C98FhflrCm330ltKt+smMQkqSyzRM
D81sSiDyb7XdDoEI5lKZ49XR2bWxH618sr4abMnlY0Jr6xBq8Yg1FchSXzKWK/m3HivzfXgR/zqJ
tmaYkw2cqDwjSY5OeNBlVtqKmSGwJdOWuMDNVJJhZEjQOoSn9jIOtDpsnvcL4groBtAttL+6CNYF
hFbr31xPx5YqtOk/OMvAQH3zzbkQ/e7MjouaPuR+5IXpBq4VPN54CPJMQhy3CcW05JduXmoMNcKF
/34FgSlckBaL3RTdZ/V67znK/uLZLH/eV5waEGaoM9z9y44aCbEgNHiVf0NMTRi1tm3Z1RouVxf/
LX7wbhaMLI+sIQqppLKKrCXK+zePIYlmGiwIg+LE5VPagXPNL1aYgZctyAjWogmsAMGbn7lXDexb
Mzx7wpz1lNbORvc+esfMBh8OWVwQpe+8eHk3s4mDj+SR9wc+23qDkkPg7AX5PEySO4blbFd8Tkbm
ai6bRaECsk0L6bE5kqSd7TIFb55YtVsHpBDOdP8uizGrNh95T0ur7jJJfa5k6hb4fy3ZlhJDymc9
vhjRpXJgEDHaVFILc19r9d5qWXf+4d0Uv4ye6n9C4SS9Gs5se8py3levDk9J9y0ldpi9h5VdwO3V
br1M39Ic7Pwo+WqTCoeYsYvchraGRdHweI6HmSYZUtL5CcgN2G4uUn94eY+DG5MH243SzEYisAF7
9O1Rwbe++e0goD6jiiRRaQK4hc36n6foEbkRxlR+nyYG9OBKvpnm6OvyCwyxwzIkOyd4YHL6Opyl
u3ruXFS+B2fjVq8bgmcFnMByxUPcaYgVKSVnNgS3d3neUVc8M5CDKMJufSry2voku4fhMqUIMONV
GnJ3+s9K4qPVN6HhCKrNyS78XvfQfg9sZbz9kgQLxzGaOQ8X3w33sbW6bxGic5yHpgA5LilCAaAj
M+ohxzT4ZRLIkxCDo32iChxOiYImU1jY/4pCBe75ATTXJIey30Nx07KYIeIBbGHi3S1u2KLlu1Sy
amJFQip2lOorxvy8Xdf7yw30GkIBSuUCVK5TmUkp8pHqcmPlmN1iJrJRWyPi/uGLxRRapul/p4sy
Y5kx54Z7+cc0LYtlN2GW/jPkNidg+x+7HhK7OfTxwEJ8M2BEpM/EB+Uci6Ip8DHHQtHx/lavkVH9
qzuiSeLbQOHW1AxPi/8B/QTIjLQRizo3HL9SwtDRMYSyAaCoh7EuXuj1Y02z9OXfz5zIEvo5iHS/
8uofRK/JzsFrilB0dJnu5k4Qcr7MpYY8Uk6LW+eRD3yf/rzZdL9Cp1RtZYTb7ocbjpJXIDTqP/1G
SE9w3dZYx2bx/ZvHcQDfGugBJ82B3EsPfbOa9ylBsmsH9CVs54fYYR4i451Z830/TI7zbKlTjbY1
w37zWU+ndIgg/sdim6n8Geowo2dFsAG8X4Esilf7Ap8Dh96KWp0A/mh7gJiiAabuhvT7Vt/rH3EP
3d2WdnbtTWIe1aaLqG33vty0QBVd1tfoHZ8WnXCzxbqJG7Z0hO1bi/YDBEzMDUX9tWO2U/Y3Lv6q
zxRo54iNA236TCV6aKxIOybvL2w4Pwxv0Gj8Ah8vxbn+RWCJAAwxM5qxmYnp+4MKpHm3N6Gyqe95
NP5UzyHsuUx/7pS4+yFRvi1x+AJJaYv3mLTJiJxiD75rkl18G4eb+wt+6wOMTpnY+hY972BFrwFL
v6An1oSulQPBCn2NnNRRFEC2LoW4uqYYVmQH4hCcGyLmg/zli02mTlVUL2MRfVjm9bjsmiaKUk0W
EShE24cKOau5YRfj5LPOiszbIhQ7DFWSQz25BRhCkyj0xNUlSGc9sfC3oKSvoRcPBuk35lnIqGJE
yoGLBcWkqbKbj+PDJZMvRPNXllFkJ2CaCDD5HXx6aNbnkq+QauHQOnv31mHoIXd8wsDo+2AmfCn+
t2JyzODZF6h4/j4FVN0ZhLQQzRd1GdVG8CwjKR5RV/ij+fi8N9O+tEz5wFS0PleNdBZOGDYkqpGX
6lZSgOoY4htJDTmCYS5lkr1K2AXEm01VGOijrmednLViIzieaFfqmeXXFb+KObIo5R8BGzeH/u3U
TN4SEz3TpVRjzwjdi+XeU1J12TvxmI6u1lWr/B7t5H9yAzH2M/l5LV0S/y7wbUoHRABH6J6ZumVu
H3caifKf0UlgzKyTmv6yIDOxw4yyhh31yEVVoCthi5ntJQ6TGsKaqqVw9O9mGDaW5xDAB5qtar08
WuNv+nci0R0O4NQX05tZbRLEBwODt92Ps7LN3adAMsM5TuAabIRu+3ujVxS2SC6WNknfPzSo5/oI
fug4n2ScJ2Qng87kH/JP1///pe4weKiDGGb3yn7NzXxXet+xOeOtUhDTj9+R/AbDWx5/T9TgIPva
hbJjwvcyw0LkUaJoO/K8aANlSaAS1Kw4gbkdesaDgQFZd2ba1lie1OdgJkyDd4GuwmO5UI7sP2og
fJjpFD9243W8zjZhqKjf7toVRPcyhsB2yFhFeTwenebmsVEQe4qGr08QGO84CHOd/S6cYM1x8wK+
nOX1d7TJzJ4PrrC5Y3fda29A4Dbr95nsQKQrKRKMG6NCsAC0j7/Hwu048YPw1Qnl5qYWqfZXatHc
AFo4k/kvcEW2XbvEsBhYG3698FNXcgVmMI/2sDLF/ayr+D7t5HuD+VtHhmyo63vGH8WBDPBrhnJR
YOXI/7p4IgkdpuRfoTK+5eJW67Xt1roiPfljjT/2uMuO/qebw7yvmbwxhN215F1YLRSIiiFS0wBY
Vippt4ZkkfCAV6EaVr3sHsQT0Z4iEm1RPZl1rfaSzrRwggZ0lC9Mm54zuDSXjU4aU4ER2QUyqRBg
TiHkcxHPCeYmmWc04/zH7dGUjEy/Mt0aWg0qDtnpy6VY2eqN2lGuiAmIAdTMnzp1Zz/vyUCz04Jd
ukbqe8X6ebZZjfrI5lDHtN63D9++Y3hdIYuusEAIS154aBUavYdog9uxMEiu5BCasugmUshXwJHR
HXHtT2q00s+So30OYQokugKP0nrIT9q23x2NM9DeQ087D2cOVTJ/Qp5HaATMorAkez6EC1Ii+Jvp
K5Lxb8x3OJrojcaYbOnV0R+wLKG+n9nlHZkN9ggwRW0BO10YWyeFwJ/+3iPI82i2Ogf1Vku9mQfL
QbwX/BWi6h9CglKgAyKUpSD4VLWyAaC8xqG7Ut+DIIQ2hErP6V0J8FxKY+/Z1Db4w0Lf0s8WeoJv
hWUyptiBH35NxciTxlUXhoBSCgTvHztA3SO+/pfK/thIHOG+bI0Pz5V442hae2KRClimQ28puOoe
2QPTqpaWp2bT3inwAYcMAq0r9D51oxuoN7dKzxH0oiD1fbCMDdFiJrrpxtbP2CIZZy8QY4bSSO49
H7ZQDCBy0yPQ286fJtNHFGCr8yQiQvtsV9Wrt6iSJUV2wgxrvdWor2ilGnQN6PFFAF6yNJGAY1DK
1rQN5l4Fq7nZaOniASFgBkI+x/b7K1zLbxw2as+lFsff52aJqFpwHSiuO3Lb899KMKXObVct8/X/
7L2oRXiK8Mb/RoLa6STj7PSkpzpiRRs44wTTxcRlGlWpMrR3SsnFZ5LXMDzRiz9aIajTwea90QPS
6vLSByFBDf0iEcrQz31a+mRAunmoPTH6riYFz/kGHx7cmWmd3IlPoig/QRczTJu2ycVbh+4k8OUZ
AJ7H/lnQjWfhb86hN39Bt8oCfFi40627FEO5azRsl8x4QF+/VDkezqLYQeaBBTVQFtHX5IQjy5wT
U8pYjIoIwlu4mcoyj58ogX0lpy26dDKLEUpypZcQiSFQ8Ig3u9GhtvqyvVGnQxBXgtlV1hXY6nVO
AqZdxqppq1wvLUSBqesFVm8wXBKjt+HifaM35Q6Dh9+zYOJXmIt2pTzIW9CqTj4HqmfP7Mvcw9cc
t8iTtS7sLHjrqFujLX4oxfSW3ECpIB6skLp9sa10GqpxweI30CQ3DQZNfwPbW/pLXtKHpPRurT3O
d4PEPP+zUO2+/bKFm8x2P+gOfEGhfupGptzSW0Nq+nbVR9FKiL/H/E20uVFttVLwQAC8tM2/2YFb
u7NX43lXncia/P6vK5urbr0BfpQFjYP683SK2S66utUdzHWhm9vhCOgfvIeCQUbAIBQ2spXKVjEl
R3w360ioqE43aCoAHSNoj+7X4LhGjDOB2/D//j7Qwb/lg89lNJNiSWjt6civBJhXGDswIzh/39n6
Is1WS1tUVum5wslpzNkrJf0aFAnnyEqoOlGDZN1FvnsylKmMMvXR3G2bAZ7PG4YuY6qpJ7v5LJfY
bSqoqIqHOf+UNmLvhu57tdAXnh1McuyURRuFY9jx1Qoz/QGgPfY36cjz1OTLES2LnA2d30Z7LlpB
eQpXWcfNsnI/9juBP91lPUUEG9plSGVpzGHKpprAakGwghZ0MtuKxMmf8HK0y0Ly6WwrvcJplZsG
oSHIWNFiYSBm0Dvm4EgjPGuCLvD8+bn/6thRIqtZQv4uP8JcKxrpjT4ttjMGa+jHGN3U9MPhOreE
LMCScCNC0UTGAu9zwJ/13LY5qBO1TZsF2+lG+SJaewnqG2OjSreUeWeCt8DjbEuMApxqP8+G0JTC
E4CytbcZp+vq0vYaFNuIfveaf0fsPuSb+9oArRO9tUK64VKqKTmAUnAgAx5Qu21RJnJ5HK6EhA0Z
py/6jgKFDhbMpsosl65F20AUPYjB3VF39OZra3yWA9s0/Qo4DZvfyJEo8BiPy5skHZfGm6iOpDqn
l9vvpyMJm7uIKxljhhu7O89OAS58B68r4T81DSzRF9kOXgUbl9cDouSJ6AgbtW/OTJe0lkAwdxot
rlwj4HC1pgxUfZIP/eeLmtvXk5eNm1vxBVfhfjxa22vXezRTJ9VwdI2Xb80OkB05KLf/tjkWvWET
/59rP9YXJJcpZ7Q3Qaadf2c7VSuphEydch2pB49uDXwcsSpMly2K9j9UfqOtEp3FpO43AJK0z3VP
3otx7M+5T3W2fVMi/eFGtZD8Iq5uFZ9LdIH+tek/5jc5iXLWZ768FnQ4A4eyEaHpaf1VlI54RPpm
Xtc663vbMu9byxyUlNiUu79RnH9cKVvu+uPm7tqwK/fU48Yt5OYxpECsV0FsDLHKicrMJ1LxvTmB
xcPiSfQl6MdRFPzTi6di1Uh6skISS+roHF0EvkhCqaeNrZ1bWo4c0cTcSjjfLm4IG8sTTgqgw++S
AaFKsf5u2mhCfbxBISgZO3xCvGM6oBvg/iVf4IrpkADYIaGPwQVGWI8U0Ms223hHjQqEv0Zg27E7
OGcCvM1SiilbbLn3dxpBhczUoXFk6TQ/4MpkjtL6UquEq3WFNi2hByW5ySYgnPKMA4BLhxPK/Rfn
7FGAuhPrgvffSOT15QsPBJmraarP+7sOG0oiLOV3nug7nUoJIr2Ly1DI5pmW3mW1MftU+wwGjZKu
uAFRBDcEKETG6nc3FElMMKYZ+YwX+EBsPkOsgU6005QWooeToo56/FCm31F3dZTWftDclk5rtpJb
8Pir9ZHK0OIFN+VIEyEqCfSjB18KUFRt3uKGhE9wHrxSl6peyYfgxUhkORhcjE6Xqamc/BisHW7R
Y2UBG2gMBqT8VVjL1jEGw7GXf9WGxSruZt32ELfL25C7iHRLiItwja9/RmY0KV/V+FPpprNMUokl
xv6FwtIskE1jaqJk+x272gakNCsgp/dbJapT+6ZVX8ylbc2yt1mjPRcqjUC1XhwSXowfAhuLd7a7
2h7o79jnL6BY82iigRnfLHX2dlLxCcftMJhrcC2fJMNGzPEWEylL67FlaLtovzDQPvYmHBkdz0XG
fVWz+I4DzAg1hRLfTUCAh6DYnSAGAdU9nqd9+HS0bpxq0frq+NXMVkv5T/VMQBb7ZpqgZCCWiukF
rKkfWppQ6OtaiOE8DrIOyrSh9kfQfXel2z4mRFLK3m2tPTmoqnoDr01IegVDIk5sLujvXVg8l/rI
0r5VI9kQ4MaNgGdou9EstApI6j6dXbBauc/AXss4Jy0+WSdN/707+kaWOFTNis5PSNC7K0irnpYi
/ttZxeq8NMCcuPPuzza38fZ1hucihMgp7b2MUmSXuuEXCz3a0uTk5NytXTcco2v/aOdq7eKptUJU
MoeR7cDPmUQ0AbibiGA+rUf0FMKSL/+fSrRftpIA19Ev7hEgwtxAUN+NB+jgZa14M4aNH5wDj6Cw
DulDzp43t/GmUfTQZ+HXkRehjetFCzuM0paO14znVg7DeyJp1Rbg3lAGxiZQo8g5PjdVS3qrMktd
p5uRwTg1e7/kW0QZRQyOo7sPHiX+UriAVRVjdMZ2HyQV0DMfC2BaQjYNtIB4GWGlq4QutWClrITt
bAeJu49rg2lep0jWjyaX8guGiUZWwfZCW9OMZbbw5jjMvTImZ6VfNU/8Y79iLVtCMe0VdqcFHOsd
uC/9IFgVTQd+gLqbf0IWqQy05tA1Sk9KoE44qmSFSuk8bHFJde2TQHkV1cyGJ9dWMaW4vcl27Lw6
KiMdhA3/Fn9PkUQJebE4c634uVdj6wYo9SvaTda7agKDxV3kpAqfOAYOfJ57U65wHkQ50dosQeJX
Ihc8k7Y3LcMLPidpKKzeQx7aa2V9KE1BWzE0kPrkZoTSw9Csmhzaa5hZ9FJ05R+BzSGJK4m3NeWi
xcJCbbQUQkYmordhf54WWEHFtLvTGbhiIOxYJRd/fGSCrLKKvms9eu2HULVldxzbW8Q17frUl4RA
qusaAwnhDvkh/BVE+Q1P/Pyhb7ownTu1Wp8ult72ih5WYFrmwcRD6ffqJoEgTyr4WHAXtqLXIquj
EVRC9HnYodxY+pmVvzv+ub39nVA8v5gS1/FYs/qzLMeXstSQ30hRggC/DVRr4iHaMQkvYkpEnKfL
Xni8S1aEdJo752phFdwPrTafhmTEdiAdYRUBz1wvcJedbWm/v5A2rLg1dNV8FKbCtYfF0RLE/hKF
cK5MAzcfxsuXIoumqJ+QWxMeWeJrJutgtKX0qdHDPSkFCwsPjggUOEJmLiMl0nwTDJQ+NqS4uH8K
kSA1+05hjhciz7v7UEKyaItuRnCCrlgQjOd9Dz+9b2efMZ/jxwx1/BgcHoTO/vkuJRwxtUZ6f8bU
4EGRaqRGHh0hTtYSUK4otat/HT6QTDIcXMfCRI5bj+uKGw8VaaUjZ+skip5d1jk6pjg1piGtuwFY
lQpYPv1NJaSN6YYfVed7O9p1LqG9dKwbAwat4NOdtONa6oqG02QE51OJ5s17zcMTzHENcronMSRE
XkAL1vU10XTilxEomnwBYVl5M7O8+GAkg1su1zNg6ZwlV7OzyemH6AVt5lH96Ft9y7ArJTZMLIrT
9MiVZI/T38/X3bUf7U/r4pNnxzlmx1J+0iAwZW58/MbcT2U3nC6m2ME6DIzRIY216Ek5q0EJd9/P
U8vVV9XEK9V4xDDtgQqoZ7Z08pDkZCaTJs6Mxn/SrsdnUj0LSA6/T9lV7jMzOTUhEfVaiWRcQtic
fI7DNR45tqC3iB4FinYGLN0XlJIkccor77n4hLGwXE2NtmlHq5gY3N8PHI2ZRYo08USqPcb6lAPg
GFCpS4zhoDW1XTD/bqf2/gvtEYjfkc1SU4xwQ/rZKw8Tn8jezGHkqowlOLNh2UTZNsj54SCTCCYO
SBp+gKG0wo8450eHYBU2YWA8zwNwh5/Hu24zubmsnmzkA9Ydh7vF0ct0Ocfa+oz7idCJr0gNk0mr
mKJgrJNDlMM++TMrrfzR5tGDkdcmVmPUem0eesjJTiedAHuYUwJbn0cDEmI1RX2U66hqCqB9QbMi
tO+qpdBGVo+yalsHRcgn/+74CxTboBDYXxeXOzYEjXMJjPv9D3N+rykaZdAPGHtnh0jSsAx6fWmd
N2UFD/NDUQrOFzfGPt87QJWK20Zypa+SfO/vcKK/74Ltxo0duX/6RzVPf9ynvarM3y3wdBcFMq4f
m0mMgJogW8+cIJYvlTX45ef6j2bpCnr9aTLygk0YHQfNa3Q3GICojH7EWiDy/UChDPQx+iJFBfBt
V40maFMAYXDXnSRB4jc3zZarBMZ2v0rVKVtcvEjhuOqHndYmPrVJAIPJNYtyZyYJ2uFyvQxFzctO
7Lbu7pwTZygReL0D6uoNTrvE9SR7csrc/0ygJhFD7loMxQijM/0pMlzrDwUCVsYESsrqspmLXVBn
hi+SkzlW+MOobn+v/3XshQoIJwLVgG2OoL2+kifz/4BiVn2DjthcXraAh9A/bzc93uZspFz5NRHZ
kebWu17p1vqYGHVAhk9FN6wSG3Uf9V32Sh7zgcsy098S5rgF/6KZvVTGJ7cMzDq3zRvJ1br9vpcO
IplffkuYDEPl5uNUpBSmMKcS+vZRMzem7aaqqE6v3ps1r+lnL4SbTDv0e0ZBaxjf716r9gpYZzxg
zxfAh/f9xePlWny76DmTDTvSUpJ0aHcKVu4TeFLAJ8m9GWb5ut/63SXRDIMBZmonQcfmyisIQGOx
1KEYqQlUcttjr8axn4fQlkwF8yuK2PEslHejUuSV9JjQYSWlRHqB+npfV0O00YJmCMmX0cray/oX
KIHk/9LGlOPHN67dqTeOI7HeXcaUpUzvxRDpwzDpkvSTatR+zMx7nEQVNKbrLrifuFtEsdb3kpb0
1+lNHTyk3R2PNy5fv4a145zl3feub4agNilWS8Foh7Bq/0fr7u9JSqLF2FFfDPFv0youfgdAytON
ECyjK2DJQzvh3ifG1186RWIlhFa04twNtUeIpbTljhdwManq9spvQdDP+tRdiDM2yu+p82Y2mKUq
MPtiMxkK6o4nmwknSZUUDUcJwAteFe5BAAXVC5/vuDdCfGhc2RK97dqWayyFhi7Bpmz8+d3p6C6G
Ff/AxYwvmr+pMKLDBrXoFBjrn+rMp50eYqbZH5IOmXSb2dizW4bU62Vl6xE5EQLDRx2QnX/1pnSR
/8j2ILhHJSVkVT6/0JDDF3TENtK1xd1QvX0sRuSRWjsQ5xL4m9YuCGSgo9crlMVsEiCT71pPP9o+
XrKQP/mPtpU9aUbiJwQEpaCle4clfkNCrbxr7NtBzTFjWth4cP4frWvGrLhBnlTvFV5sQ4ixKQ5s
FMfqYS3GpR61jhJC/yT5TNEEwMtEK3M0e1oZOH6V+0lrjVOsf6ASmgCp62o2GqJoZSWSMWTrjxiT
9TSImgeoEls2RsFanz1VYHhtZxzM9MsQ+8Uh65bc/nAqZK6bAFjLg3R/LFQJQ9KfMl/56jwscomI
nTQRy+ZpYgfFBo8794I52xiWNh88Yyp2NIUB2dYvcPazoGNMSLRxwjhXA6xuojLSfUpq8bUQnQ8z
FyL3ZCKyLhWajnEAcsCE5+P2VPONgbTabdk0MAfLCec1IYTyacWrL2LCvIVUKwow61lt4szucqey
WnigcIesZjgdI55foM66YNMTHSOEZN2XHKyRbktUTI9u0Su9VdKLco96TA7x34+kppKVLTU5Otfw
fSUO2PGjAPhyBv2YI/wbDpFclSraMJPMTVYvtG848mrsD0onJMqWIDzjE0mgElrdxmGoSVYLR7wh
A7ssZHGq+Op3DZkl43d2SSZc8pXQlpKhURk87ha3m+Cak25g0IqsK9TzEvE8Ea22yzEsBqyT89IW
v8vZJBO4rmma0Qvl0W8QarAGsT5Tw8Ehg2p+ZmfcZFtShx1VwOdpxUrCDhqDHvWuXYgcmODNNJyT
UxYy//4IjjekvO/lUKfosL8+pIGwQ5e1UVkysX/YNZNakufN4brjg7oxPKNyDlZQZtkVNpx30AOF
STRsjp+sA4BudgrBLm8HrbtA7QqbUAtt7I0qG+QLivSUK6KgITulJjkFLJzwdU67NciUf9r2Erpm
zttZ2Tn/vwQCRAWQcF1B39mdhlgXh6UiUCJ9LxjNvoW0npAEAjZVLteGltOD6Y2t+OBzzRVKhAUG
dk2utS4zJYQQ1/truNKrtKZRT52k5k21yh9wnbGvpAeSKbraSjI7Msd0DxI4Kj6SyBFj0F33lDv0
vibW1UCIZ4aE0qiouSE1oS6wjOXf+GVZ1jxQxhJQ16BAbAm3y6MpL8UXrCMBqjSg50PVdn6qEcD4
gPjmRJyLwzi0ngKZclkPZxUlC07pt+l2o+9yrziUTxix8t808PVsbAJQ2szd3ySUkxtW/1RbYSCE
QQ/WXG7xvsm7mv9ULfY0ZVy0Xz1fVzqX+fuf0KBi9sJ4WJuoDOkI/GEEQX87/+Ombn8Q+Ujz5z3D
DEQJf4P7Yi/54DshfR3IPQn47FNESwjkRkKHtakjwQkM+x0BkFogWzPdnt9y0fbxV2jXAbEyux4/
MS2jI74+dpWUgnA7wHk8xzH+zxQTXx0BKsJ8pkt9pkFsCOQFYhoswXfqQCpWBXcrYh4J4IrUJiei
2LjLkw1zb17TBjlflNn0QUs8p4rjwVOQAW8qGXcCCrlcrYnyzh2VNL8HyNisCSoT0g2wtj/sFwY/
gEzLGHtIkLA01Vs7wRqgQt35bPnoGEYeGjD7CSkhJufSxXZ1YcA93zLM2kNjHQD21nBsRoHmAcxC
m33qdB7gF1/YKNZjDadSb1ocjdBZXodY4kcjOIenpSR22YG71nbB22WH8L90AyLZvsyNQAjsXIZH
O1Mw8ynUK4nLnFWc5F3bc8W/6217rnsld10KV7Jn9Sceo3XqVSUSj4qmAkythQb8Gb2NJIDlJJCb
jw0hXNyEHMxVS196hcrmQSTe3F34aw7VyOcGL9pWu4oXyCkMjtoku2EX12UatgwZyXHDperud03w
qiljCjVKNKNWwvqWnhBsx0c/3tKZ7ok91R20LvdRpPnfeMF6x7acU7Ud1wPmIFGqzJm1FSUPIfl6
+HCq/Pb2mMonj4Scwl6SxHmFt7ZE1TqafwuWky76Tji1c6z6BuZgJwSQtAUIQLL+FYblRRIvEkxX
ahzZOMe/sHXQ7iqzoFQ3MI/hXnZDg7PavuUbOLLbAEMsqg47xQXQ2NLcIW63H3vCknhgS3ycywC0
Xyqsg+KYzHa/n580kD/90P9GCOlcN0PxMrur9Y9VKT7AMCaUz40qFNNjWKctMH5DTsaPUBaLxjzU
nd4BiNRW7mLYAiwzvsQfVfMaOVXlOWRhrk8z+7TKNm/5jFlGxm7L1O6PItDUxQqDflJfRiVIp9Zx
Y1nVdqGbuvmwwsfCXb7sNqYpOsChDk5+X/VFqK/HWVdgWGUgu+JIJ7D8QDAQmWtsmKmi/AaZcJnb
lOseoZ1LNMGJh5dXjv5VufRWak1EqYqo9YDYnDr1d++4c9y0SzQX7Bsi2ddOCeTNMrJhkKglaFBX
bzq5s2pFELNYjR99caeFuJOZ7QD0YEcPF+Nu7VJnP0lXl0x/tj6JlzInlmjJeNWTIMGfJUqVepGz
GAchkAWAn1jKj8sOkR30b73nA+OU9mpf/4XL/frAut0KB/HGmk0Pt/tDQzrYPg635YHx9ToUPMqv
gNB7Vsp9CHGellOuPX6X/D3MLLA+Y4hCPyzry67HP3JKMpfwZP167uaKcmNZTvXwyIX0Oh+TJGO/
ZEgiQ+ZXMqzC5BmmUtYDg5NS7cPafmf8bd6Ij4RGb3QZrXrBCWbrEMeZsomnX1x7pTVb8t+h+xSp
Rndy4t7wH9ULBE9FwaoWNhpwxEnHdO7aDcltheRuGwuENbRHnYiGcjmgLxMSV/3D7mXnKGTNvcyi
GloVdXZJbKnj80wN7kiLCjzV0TuZnc3vnqfJyzF7/s03xu1/1zU15IWMcL1QOQz5OAu8EtWo/Xqp
/Fi7ZUD5Fz2gmCMUivfclGDXiyk9IsHgWaBFklRuyfBSAWaoCS1/NPP+ma8wL6mkZTot96ISZrn8
/wsMV4MhO5xMzhqIjt5qAUhCxOSkZVCv29sHbZ084m2h4W5mfftdDOeIqYHV6VXaJOfZKAS7kCQf
8ghzfx/yXxlNsGgWqUVIWtLX2W/LGwQF1PCIiS4GLbCmGirdP8i2PHK91AUUB/5SHUpogorEAHXy
oJpT5xabQXnjgj/0i2a4A/NYsODArbOVA0UFIj1BgmwUZf0+mX95SUp7jCD/+PB9RY5DuQAONAtt
EpXXbEATpzPIKce3XQDiC4mJth83T0FA2U91wdijy2MyZaZjJ6dYKqvvOq7iKHWHUCzozKZo7GgM
md7FvqhhtI4ooWkyA5/r1mSxZmYo2tKmdWwONCVFZ/XxSUAcSDMZ8YUNMZCdu5sYSn+HC+hVF51E
x6p3LsBcfQieEcRPbpKXqzAo6vhEUkZ+uAumW2f2wsyojtBab/mFNg8sqlCp7AvxiLafyga22nx4
EPrun0Xh1TAIffAJccSZgbZVCCGVNXeBq0Yltj5EcBttScE7Rbi/MlbLeK3vVGjNEwyPCuK8kG0X
YMFW/cDC+fYhRpy6IsGlFBW1hE65f1KG83PbA2mZLuBlzrfakOM7TD7fHsBFhQn+LlYxIO40VFMu
PbuUBbg6+rABueU8qrvM58ohjVwj5ygCZhFeDuup8ss9qKb6G4JyjLFD126e5z8ovDvXV8HzOlpY
6JSFSkLQHWgBkYkEpKIz039vRRabq6Z0DPhvmeHLzeQvx3iC6tf22KnSB1F14Kz7c0rqWJqKdd8X
9hf8l0Ilu+Zz1MFOJcJKaibPtwkYsShIs1EVudI8jWEbvEL3sgM0VLrXHkpFIGFRavcBqCyFhogC
hGVzOaHPNpme7frAlwq4RMoUoeq3C+TAauReBu917amAJV3SAfT4yFW4fU1TBKC44nhgAUAr/0JI
ghl50N7aM15k5tqn7MHqh4JCP9UBa38o9idhqukR/xWSKdO+iXvrgBZ/OjyEx3BlIv03pA9Mp5d4
dVGySJKptn0UaG0DmUXqsgUGEz4gfNIT8Yco9yg/6qVJK9qEf3e/q9zT0LixIY7muZ8cs4cIOeeQ
osQJ8UNHTJwo07ZejVzlvllUX+pnemBZCZ4fPi6mS56K0mFNrsG2NzdjzPskrRG+X6MELromyWir
pjq3AEDBHW9+/v/mqrcXwBpHE4sSxgO7y/k8iCMLo7dwQ6QtmNy8ZJ3xK7HijGe2htvDWE0jl+EY
H7rmK7Bk9oSNSaxRTMYt8gpoeEkZzXCaZVKosKP2j6fDw4Cg4jdwxgK6XI/AjOHEo5uLTiToPpjW
d5XVXo46VKNOW/VIhKCVNAoISH/76JghzHNbp5kRMNPHdOjMICwPXT3zBOM7ErcT/f3zXZbHA38/
8uekpuu3Aus7m4l3VSxUZrmWX34T1o65XNe2K05hLxkVOQbSfdp9oZcsupcB8Pm1gif5ahJyeeR4
h/msJu3DAtE4qr6d186IbFsiQDw0FUWw0G57/rPaDIC/z6RFI3loyAkdLZWmaQCziZRlPay+LLK8
HJ+6ghpEGLmkj/P+/wIvtwnW8/9YPMnJWuiUAbwB68mAfquF5D7vtzFF1b+9Rawp/g+KvSbkM1w/
ETmAQjw5GaCApRfP1hrFskq65Ut75xMLV1uJy8hyKb+O5b7KQ6Cd4jus8hqIEQM9gkI41wq1vTp/
+FF6TT7C/JEW3xvyVEMk9qV8WeN/tG4edE5bqE3HsusidUogjxbsv7RHFp+RjZUQvu9a8aPSCBTU
D0KbrIBlf0EqsMiZGrHrsFLyvz9iBiWA0OMQzpUrKYh8rIWwTAXsa+AjoKJcgdR+mcBlVZFldK9A
KuWaB9d36WT5rhQXjqeYzq9rbZ27FcYGCRcv8zeK1OP5GSjD82kVCkN8zCBXbv/mQN9no27/Np9E
ZPe+YKwaWDqG5G9+Q4pF0c0i2OVsbHNRuMlf0S3D0acW79TNa2VZHxecxozIesGN5uJcCX6d3sis
15X4CWPwgrZP9RE3z9MfuROJCiqR27FDemcfblLHyig6H8njjqmn1D4R8IeCZ4AesKG2d6G794Y6
3MTSYLBaUHKY4Wpb3dSQORSSNNbzgZtitwsJHCJv3uwZdbXAQRIMyk4ivVDPtjQcGnqJFs40PjL6
bcpZRyuYyLSbvscT04uZpBIkuERv7UdHSh1g8fI6g5ZQgWRd0nPypXQqLfHvAHL5ozLw2phrtat5
ykrvnI08QpylPq6AbKCu9YEHtVwCEjtOHeRlKEW50wFjth4imRFt8XV0GKyC180P08pJPkLePoxj
8BQCAC70240sfOjoT55g0zxbcbJ2t0Cda0xW8mr3PJ5MxvZeLp48rLC+Z+NOXVQcjcXxoSU1ANk2
5ZTqRO8BeDuWM61UpB9QhHaEkjNazfL0tivExKy2rPfkRK7Gbly6GkZIemmMy9MtOS8jBdOtmvm7
ciKhuYp33KYgAHByw9GI4yfnZ6GUzRNitRj/QXcPyv2sZCGucjzGLPUMOyEvkyatUdYTuVArDYEc
8fUuFyynOzAcM3zOITXdQEEuZ1np3zP6bvzdd1eSyFQZQHh9gtG6V4JLbGeXPSLmtBR5WE17RVFo
BhFRs61pAXAfmpGUHANgmTXwOLpGJ4oxNBf8w6MPatFzAHWKYHwBp92kKJz9CEeuMBCHhaK2b4oZ
hCL6HWNVqIn5dDC2gmcpCFbs+OQiDe4skp4asFmS56jMt4osFLXqXQafckrw1V5zPWIlFK1NOwC6
Or6laxQLGiiMInnWb9pTtUEu9lN2bBWXuRkjteJUrTw+8Lqnd/h9g++mdzrD/YoLSsaChAtyxI4Y
mmhiJVmE4KoNAbHNmY032YjZkQFUnyOqQRLN4k76347zi2F3W70dFHC9xhQtEdoeYqXoIJFz4YJR
kXsaM5v5PIES6F7BbWN9sqJXotGwZvzx4JvdHayAmZEkNNeQOgxolmuW1+PIeZhTrrNJo6+aUSqN
DtDQLcrdRty0fvvWljWO9TTIyrvej83Ma84zRW6yKdEUWi/GCurFqop4MMrEmhGOvXcPAkDLNy8v
f4JCpXHsuK4F5EEXsFI3yyA8+PB9HKvZVPyEJcBWUxqi0wRhLfSoskrCxfK+xMOMLdkaeAvs2D4Y
qmWrzzsVZSbtJn86FfYz+CspidR7fW6azseYZpMLb5NqJ7xrcmR+itN+6KCOc43MIINeBS5R96wy
Vy328Bj2pLJOc5C0Cm9woi8u2SMDyg17lfGYK9NW8mQFz/SECA4UadLG0lGNWG/U1FkwNFZsNc5+
W47PXiNsFTvEwZqarGAx03bd0iOhD1EU27hMya/6j33XLsciWVVXAGjNxqaxWJShwvfqvH07QqIt
I7JAkkKAE7rcAi59kpjGxXJcfsM96GXssRxscrFUMRARAInyNonkSSVlFsAHI04rzBG0eMPN3Ygf
dovqzcX8KPB7eTYW6D/5MwiFuRyihLmKj3a6sLwK5o61TYkNwoOjm4O2m2W/oWYZCFGE5EK4yWEL
J5/1TfegEef5Zso68hat7DpyBuc/tN9bS0WZXKmdeHVlXEvrj+4QzMpae9jnZlctJyX6FCOR2LIh
Azso2GsfkqgOmCsxKG/jDYRcksLd9WiD1SCUyiA74CF+gFf7taMU6lFKt+7+aiOGHAgkW2bHODv7
ZKD++Yu2dhx0bodparwtbXXb+SnzhqSjm/nWpklmpceTZzFlFMeuz8yY4GdBdH1TFxufD1aeNa4Q
W9ov/y+7a4TP0Opn/BzniTquvo+0YHLWMy7dhMf7pifu8qo4TcA6d/nPDMzj2F4btfM4WY9SoXp3
t9LHBt4VUqIuBN5G8/8OsdFlWpgPVqiuhYpjceXmTrndnxtKF6iKPawuXDSWKhPlDKSjaTWq0chW
vnIZ7slsF+xJmU3ydYU2zv2OuV0K1f3mDX4poHXpZqaJ8NdIjTGW97/N8vQX6y1ldpgT9amT+2CU
JT6K9K75N28aHqC4bPZa04J+7wEDBAiK3tcWaEBocVcTwfooMiHc4bfWi50lPGAVSYQhmp65k4gU
NAW3+f//Dl966a9qZ2w2M4yLBxqnZRSY/+GFBKoDZzE/HSh5IfzRXCj/kOXETeCK6tuJ1ShIWk3c
ZnXMjMLFUsm4GJQuMDjTcIODr/sbqf1Yk1YwH7RzDSpY5nbXj3/QppaH8t5ZM8A2iEDN/olZe1RP
6/qXRnBqMvZsSoQBSQNCwEaQptMbteYB1IQ9f6BkRbcXDsqf41Hmn/oZpl/N+nyAtfp+OZbRMKT9
SpkYham4/Dbdev3pJgJB6KNLYGbEOZ3hd5jcxkyNI3xTsYI01icqBGVdk0+Y73BH9Caa73bmXxeJ
d8tSSW3bzINXpIXHUsIt7YYvAq1btWJSq5XrG1wvCOUNd/MElrpGyluJdWUc9Ea+rlIKmmKvx1sm
We7GWW5Yy1Q9g/HB0kVZXfnCbcMMT0nm+n/KETAo8CV76SJyZPheBSpzsaQzpVBZE649S7ppcO/c
8aDIzh98OOwJE33//m8kPj7q6SmaxXhEwmwmHa7XzFUD/uDzVhpaNhzQzpyC8zFeh+FolDL04Yt/
8/qU9/Ft0BLTwHFCgI6r6nqrpg5NMYgMt6tqlffQtbMlsy3E+rHAbwHD0PhaXBmRIT/N3E7gDRJl
kwxosRhm1GUroB5VWdhJboecTq1CBBHtlworPfF5JeNavsOVTfsSMwcam6eKCdL05Jeu6Jh4U9vS
591NpsX0v2l8Np9pioVFv78GIW0QpLyDb++so570gqeuLzkmNSGWG/ml7VgUEm5u3onXGDEI0WEe
gH6vS0N2z+VVeizN8b4+jxAcwwVA4iH4rtp63R+sQpideu6j+Eo1B+lASIEzb25T4+oYxzuc3Ohd
vR/KvGo7BLEI0oT47G06UiMMvjSrWxK/oOuI/DsyWWnlvlseyQVSWpQ6lmNtTCJ6TZqpagzsSNWm
HC/+95/VDtb2+551FP7aGjgSh9la52vNaKUSOKwu/9vGnUWqHVIi72P0g9IT7GdirWdSagDL/XBy
3+PmW6K7U2H5/ZRh5AqZ0x0W7vxMPhnXKxLa1SOSz6HoGt8wdhyqBRM25NFELc0wWH8ePiv/2F4/
gRe3oBiP9u4ErGUDEpNFIIlC3tE3ymPozFtIdJu25SGGoPnhvzG9HYIiI3SC5immTgMo/WJpXA9o
B1UtfjmgAyR4DEaUfrlY4Yc/pDzm7GLlEo79W/XlzZ/KIZVG5fZoug+eGvYgnihvKtCPOxuBAzH1
VyRKNCBsixQiS14fC3YUNcEPj7l1T0ku5/J6T1BiCRGAMvE6kGjLZQ+lsLbCfjNlkdYl3xlCvaaB
eiob4Pjuta5mSTCuBB6XvczJiAx3LoS+eVUUe9/ys+cNRnMak0S6rzN13m0ukUsfYmqfafZ7tNpS
6rloWfdmWHFdcD5p7uMzpxplVaFusPb5iviVxSgvG8+dE6UHUTIcG4faI0JzRCCdANgw/fv/J8df
dbB1RAOgFEBzxoKsqqm8BjHKg7NS8jN0n7VZlCEMQp1+U6uRYeFt+ckMZFyqTgs5XJnpyv9JW+WZ
GcB7CtutzXhisKl6nAdgodVIbzd7POtBE3WJ2ywkhpgQfXxRot5uR5paD2EMFtIeIb0RV6huxOR6
/oY26VxIiZEcUZfg1kcpQ++jsPHZBwL0qpvl39mNjRhjyiKqhVno58HwZpahcfKYvpxYjp7sxAWZ
PmVjW2+A37Kk0IlYnHo4SHFe0FmEi1BIa0WJ4qK48oA8NShWUid+knKSRAzegDdN0A6xQf0GHlqK
BAKo1odXXojg5hxiAhOSYqcxt/fiTliBaK1DscpgUpiTO23EeHHnVoNGXfmMtfPfqzDTGaAsAcNf
L0YS/YjdwMvsOKkB/bV1JJEse9nxm3j7RuCkdAPRGKo02dKsX8V2ehy/iPZC28D+x/mBlxOo4yVv
dwRiiletfjklxRUt15CWWiycAAIWFoSI6fCD3KhxQRt/FOKy99/nhdZDgmtwsbHq+NzJEzBkJzRh
rpvrCa7CV16vgUMKyLARBeQvQB5fp697EKOxa4SaPUflOEM4DHK95sc777GCVvL++XCpDv42/3Xd
EkCwS0DRX8kaEbQUAV3sNh16aebcwx8NGlzWh95/QZVRHbrdTtDR6h/lPwipf9VBvAtjg93ULAaj
34LW+sUQQU1nw9AvrnPbRtBrNcBjKX6vEfnX3gKEcHVR+3B+h5YH+Q7rykjW/pLbW2HwwqH1NGh4
j1i6N4doErxB42mp6j/1gkuqthCNrOfOqx/0o+ujKDKUKpHAtKpIArq2be+wTRjMVsv8ViSglGp7
snMcEFHjge0acEX4ysYw1dZjardT3wDe7+deYLGdl0QAghNmfZTnDX6ydVTT2ysnmdtb2Gpqj9PS
91noNBF5PoOs9aFBWvzfJKJDuRK9h8ItxojHU8JFuCVvDU5M/1n7/NJtLO1cXPXypaQRhrEmTNVX
5xqEkuQxV6zQiQFkg+ap+z3dz70fS4g2cXTKSjFftAilvtwLbbFfliTnD0WoKgveDKYPUdotpBCy
L+cmvbHmyBGcFGfv+Fg4FrWcbSqkTWkJmDKGvm27Kl1hHz6KG2wBIa1yMKmhuc+R4auWa6ZlHnmY
fG2dZ/JIW+9xLTKxPVsr4eFO159v0/y8bHb1OSVsSIEG5KPKx7RwAAU8+rWNk2xoieMqOAM3r9WP
l2/e/1i6KyBqbimPuMwbFmmq3kwA0oNVcnCK66+IVWc3NNv0NUATl3rOE/VMYF7p4Bo6A/rUSnpf
6evVlGHH/Q5CHFlicodfjoZnCoP1BP4I9HSC6KcZLdqSGnQ3vVSd2YGxDioPE3rXP8Z+Isl/pIh1
AmqdLSgQha+Ta/KJbkb9cIDM63ScHVTLtZ8X9NcLP+vzL/+oyZtmjdEGmS8ujWv7AnFPY2W1Fy41
IByyjoSHasyb7qzXsMFk2E8W2cKktAfY8vwkjPUHUtcRQ2fAKrnY1v6jGep2yc9hzd8geZMe+1kn
0zXEgLcNRQcLJfDJiGjG+ywbz++D1Y7LZ9ZQPyEXrZpswgscHRgcUsBaIYF6GZ9bAxVYDMoUUiYw
5gVirNR2YtfneqopLGCmqlqBlKMwKP577J50j7/8Oi7mHQt+uhyxuYb2o5QPaaNS7+w9Ye8DDDKo
zduNPUGmV/7GNf0/wOfSwKt2R+aoU4Et9spmB9PVezLNl9yVyWyn88sSrJrfRw5gV3rIgbc1qGUz
/D9iZ5SFr4Jl/TIOoSnKj5UIq0B9PQRZ9G9fD0JcVYSGuernhhfhaL6NYeNP7TKOgvmI+yH8FwoV
D1pdp0xKgrq1LJpTJx5mCy3P4+SIRoaXKuVnHtR2LBFmbEebzzidVL+CibuwC3h6OXpQ4yOmSilE
991ztADla7KIGmJKUyYaxtc0C9hQmiUORhUdUkUx5yg09lyfViT2As2J8fQ78CvLAL60dhty15rm
aBEbAHxYRaE6jaPuNqUOG+Pq0E6iK/uxawbhLEWU1u+ZZC0s+unI3op+7eTPw7k4CehURyRWaIlJ
SAQQjFNGK3+nfRvKBxgjH6zsaMc6OQqpkdSAlTs0BMWN7aFbQ8Yu+dZGhHIja2vTtR6jcUvzM+Ke
lZ7M3bZMsQYPHLWzSzyVjGZaNnOGSfDU4kMfQGFfID6c2yExuMD6OrZCgMQy7iSDnWejngsFB6c4
VXI8Do8PoFSAJ3nTAkxuMInPV3+Km7US5Xvyw70GKr9onryE+REimkU808HIdqWv/ngyrOfCZtMy
noIYwa8m5hw6BDN051pfVZWaxxemZh/Irf82q5+wJr4myizkYaOhicWP46IbzSVCwPUnkswbNxqr
3ZFa70VyvsmmWQYhlXtlkGvRfVdam5Y/A3wIMtm04K3ldJ4rA8P4l/G/8Fv+B0uAFZ8W6FGGSEsg
qdmO9z8ULgMyIL+QbLtlAY89feCt35xotZ2UrZovZUlolUHy6kASAE/HWDP+TW5fFCwz8TuP4MfD
RLjVlhHZxyTL+N9DCY4C6unr3xFtO7WSO/f3EXDybGmSpSGHPtzbpcXVoIorRQf0fnDK6Kke7drC
slz7cxvsLOIbRLGSz1Qz4hG8ypQnfYWxHyd6NaOETeksA8h1fl4IHB1b+sw6ljVYluHscDYgEKok
wjcIoNThk1TWG6PBSHLsVCm8o4YVCz1XogxBLFyb7wYpyBYiy4qlFMbVUo1bjklmh3sEdYCFq/2Z
43M3M9lR8lwBOXVIWnYClizqexw0JEDPWaidWtHCTHIWUrHvsV4iyc8QtBDrQ6TnnPcD154IsNap
WYR1YhrDtYxDsyTj7t9Pu3l3emJjjoIQaflr0MBXQuTwmAQB7WsqzteIyJ4vLM9wFAeLBlLhLu4v
tgHAEHcOW3Dbpuo8YdDVxceFfa0LdhaurJLkwYw/YDrm/Ky00PylaIpZqa6rEGafNiDqcNo/YCyQ
KKQ32+puORCkCMp4tFQdBtEMGwMIlOZRJ+k+DaZG1xaevMx9G5Ny8XWfeNJf2cvt6P9H/zJHY6y2
pNAYsOrDKOTjhOCvQVT8wOVhe4FRcxs1S+ojJnnxndeFrauH3KC/sB6USVHNjqwzNss3g4ZdZwDz
xoBErzdUty1EIBBlGBvGAab7rUWQPv62VxfpbHUyAmu+IU1679SUt2yw28OXoK4K7KgdHSwEudsz
fC2eTmdsNajk58UMT9bm5Z0QnOZZeCk2foWc8oLInNr0MPWJ1/z70HrQppNkLcOPF81Lzd1qlFoZ
gkB7LhG42/6LNFdki42vh/e93UBx5w3EpjZQps7MT1vFPQYmWatUL5g9M4R4bfBVmRH1PkZhRHOp
wFXl/xqvd0ePRzt3pYhGTR58kF0EsauhJ0LV5yqt6odjUBJl+RY6e0+ilmBH6oit8TXRQXySBmIk
sRuyYFnipN/MS/HTRUcImbhectK3xB2XcrIklRItAGS97W+zR1xZBmwdLrcaE8q9nTlaDYjtBlOz
ztoCz7dV4e6Wem9R0paSaaAczgK0GDXHJgfo3s0tvQXno81RMvGTeoc/TK0rXS6ufHc2rnALLjXs
31jY5OAO1d00KSZhUa49ud7a8chBkM33cn4XJui2fpxzU9ecUiE5V/nvEI1ireWjHujFv70g1xcq
7BbeK2ChfRjNOSIwEuxbLYxIsbFKs8lPyc4ILg32o0FIXKEfZvrNEHElTt/r8h550aerXhnwA6WZ
G04DiScHxH0zG24GZMIZtewUEFNT2hl4a6hLhf/0xv/l196qZw5SGn31nKbD0iME/3E/nb/QUOXY
g7N7mAtw6L+Zqc9FEsMkS0qbKjv5kGC/WBCL9gbRxXrouqSw4X0WescPzF0vmZfhGc4A7V6FhbMz
xyaIZUfv9Kfg73bDiLuT3i98XYp2jud9LV6LPM/JnnIhufbX+uw+oLb7hSy9WPaAG2l+o5XoJQlK
PFX2xNenQNglJ+2SWkNHedMpQ9Hfs90IVVHZxO/SdItYJ9RVq1KMlWDRqiYiy0ogiAfwJgUIZbMB
BgA0jwJLFU/PWVZYK5SJBTQsPMzQP9TD5ugO+8QGz5PTioalJhRCzN/IueptEgITn2HZV7wDXxQv
8vXwrCFU5srySs1U1AYs12/KVo3Fvxff2PU3PcyFqTjxHy3hZJwN/Dn6B47fkK0pGAolNOHKS0Br
f0SfF2D0y7HBQLT+E99JFcAClNzE3Pfk8s7VkuY1egUgnkowiTrlG5mk+y8XWAS7QfzVLyQi/9qX
XMC6XJRODrEuZxAQi32EjlG5sSE+BNm/IATmwxnnCR1DEMtI6uzIPVDf3XlQgit6lV8r3ZScVqSA
+Ij7t+BpAi1zS6ok2ccijVbyTMuiJZVtt8UcV0ke+MUYErXXXigD+mzq6AjgbfMu/J7TGPKeEZB1
EBVqMMTuojXpWxGmuYF+Hurmbj2fKH10MmiwbRCewlxvBfYGnoD7wY9hdw6NITuL+MYclg/pIS3r
q/DjzispKnBC9H3Yl+0wfPCECsOEEHmLuZTHAjDAxVYCAbj3CUiGSFvqI0DknqRvjGDJeGPv92E0
Y8+SlKQ+U0i+qPDjJAWKqAfAghzZTj3rDZyguNEEjRnBNUZ5pTaHY7T9Jqn1u340aTtmJWY+C97c
ZF9fPcuVSt3hlun5d38BGd9WQsAl4E9K8+ZJ+aLjdgrMovV0pIpTQOqFmLVfT4sTn5C6QRQCgMse
jAnCHYsrs+Gf6xurfsLImlbMJm97mlU0Ly54h/83ougRa+Mu4ZqTeSeROZXFiSZ7IRGMQ57MN8XM
l/XZ2VmR8ESRxavU/9BNqdJ5Mjtz+VMXS0JkY2DiheiWoAl0vDfeqaQAFbgIT/VyaG+c3PXGQbua
WqOvJ8y6+i+XBPoGbjTvX6RuGQFA147bv6aROLfParFnasEcs7dyyFQhpIun5sdWq+WG6e35xsma
OCqHttLpGhnkMazbR1avxyT7ALB7VULwoqZInx2nA8OhomCWzRZiKjO7Mz6qkkfr39D8K61Q3nhQ
3qphYuhDidfdvGxrcdQpCJdePUKJatozn7JHe0/YSsYUWL8nCx1X2cDn+wj5BU9MG0gF3V6d5aal
rq/5b0YIepdRkxXMxDzmeqLoLiXYFz6Zcpo0XJ6bjN7n1sOkOvfrZWgYQ6BOUVPGmWjfGzlm4UGA
oRDLhrsQjKrjA+ywi2JpqxNLuJvgp+kxEdxxxtqlBjnZHcGg/XFdEEaRbORqCpjUSgRyxJ1Uwt96
KRQbSu2nkTMuJEib89sdhw/duxufkXHt5VZGGD/fIMH5DGf/tzMWZF0N/5aTlcowpJfc8+uW1Lt0
hG4FxAiUAdveqk/Olfqu/X+U4bqnYVxqWafn/qKewTwrdA1jMBFeujHu+qDmO8zQQGKHt+xnU4qE
AyngY2u9m0AX7LMnchVTCorm7tdLWRQ0ToDk1pysZAoQNEnno7HxZCOVLSpFm3yBhEEQ7EF75Puo
Se914csovAtS8CCRvANaOiBuzMWUtnnDprGh02W9Ki6lfmdLlUwpIEl9gVCggb+/VAfYzjSxq5zp
FrjS6yJaC8fPHh4LflCJUdA2gOopQUf3TBr7F31MxWzF5BMKFkW4pdaYljXlIdbvdGfXSbPJk0A4
aHl4V7YTdADRv83gJkRKL0nKYyQz+BaG8SBwcrRXH6navGSHhfX9iaMB1ixsZ4nTs89FlLGCnDBo
OoDVVV6sCkSv7B7U4dkQGZhOtekTOBruWOq2jYpeTGojoOw2OnDJ/8J3eWjxk68Z3jm4Y8FkZRCM
hFZ+5dIXnBLRXZWwRn6/Z9x8KwNp+cXJ0AlXait9BLNxY8Zw3wPuDG/tlUIl/84Pmqyqe7e8r6Me
F6JQDWqeqww5qJRavldN9xOsxIJc0TTWequmTQLpT4gHUAyniO6ubpr++I7KLfxiEfWzxJJXshTw
PYqKNUcjl54lPBxfHFhlEI/HlleDlEb2yG3r9czP4fL4n/9NLmZ2hWIDGprpA7x3w4kfO4VBTlA6
thjRj0tSmKeG24ImS0CUaR22rWfng4yWeJl+0f3rQzvufBzjV6QB6S1mOnNGkiZ9kLogbWCe7w15
WEHiLUEUTka2ofweIIAmg6nltpEELyWpvrffDbWoCuZ3W5oqafZJu36F/fmwQooWIv2FDvmQ4TlO
vL8oVRApRpPoU1VqFHi+IjM/r2oJZaJ+sgDF1aEtA699tleQx0U8fQiQakG6weGxU1Tj34/bm2Z9
x/UMakbEjnwLlFRYaLNJE/vHwTiA5jcvlI+4tvNwXwwsXF4t9x9GFWydYTUPx1DXAovZk8pokjgp
NN9NrvFfIrpJFm6cLygxAOaigDVgMXAdwWzBiej/a60wovu6XIG/Rvs9nKSLoSmsK9SDTKp60Jik
CtYOyL84xL3l+IgRDLcJ0jtyXSuaiauXkHlgAOKvOdQf6iaVC8e6mmmXeOCV2OmGsV3aXgbJe1Jb
wVU8WcSXRX9+Y25/IHE0FVDdpGexv2vQTthiDEjon7gRApMLvR4Ve9Dhj/FzInMxvqg4lzhWM7qR
y0xcTlFe/kaOTOvDhn4kgqwuNPeZiUj+xh+sueECUIEjVsnhasrkB/6xU8lDRo+RZtnOyaj0Ndzs
eDyjCXpXsqDBxCA2Y/k1q24aJKce2x8CipF9PAf6kYqgtNp40AaaBy7Nk6irDvN5CQ9/fYf5nNlk
M/4LbXMElsy0XLrhm8NSWTzf1/WwIVupvUWsyc56shZsRc9ER9hXTY9j9dzwU5pRPFzkm1/kiDEC
hYzgPsPbFWJMKviahcGwfMAvKYeJ88DD5RSfGJsA5579rAxDtRt3zU6jD+1+GpUNVtmU6wGVQway
AH3yDcAyFHqvcBAcn5tRR6cVD2Wy+WSh3HORIV4JIah5DahzsfDJt6WvSGglFLWAVVgl9/0Dvk8S
cGqG9C9WoX8OQ4MjWDlUmRmjrIfvH9sJUzxEGovb26W/80zB9vOg5k9obJYCGGK6w9A0F3UssXKo
fF2f8/eGPj52Ujs6X9iRfFXekAtFp0tQXcIq+YlRrV72wguMeWP2ObE+O4QlnJf0v8ST8cfW3xS9
6VXYNSanokwErSPUxXswHmYg0NTKOjpBf08j8kYl7Bm4ZpQ+tqgF/V7btJYWaiTmzcHJMi8ShVP4
Wj9g+tDWBZzRueC2CwWxv8bt4HmFyDzaELZUcPGpR0TU64QoXFc/zFBe7Ly9RCpeTrSH2NyJqpyd
l/EPKP+hh34XiS3zrBQMCPDu7ihvifJgEYfsKfnfy6cTXDkakznv0O+k8OVY3WzFkpdI35wj3Mfv
zj1ySr9+K/1V3N05Hh3lW6YxwsJKdg/iq1LTbHy6dZZK9nPeUKQSDXQ/a1m0UCgIo1qAhnV8ZycD
e+yi3SgPSnq8llMrFr8T9BN4xWT1Kpy6SmCnXi+sjcRTTffQg84D2wg1QIBajCCTQfQNPU5GCR93
qrPHNeWwTGgu/ezbnrMD8SmaaPjITRwUju9z9DFjhhurQlBwyBPMA75xbxzEn0pkinfVmVeJuxr3
CYT7OjDFP7VyDQOGVsYSMPDsiSn0QJjo7vBEg2BCtWrEzKDOJskayWyTLoRc9cjvqoGhonPLA1cx
tFE1UxMgBPr+5cuSqsN/a2S/vYY2fFrZmiguNOW1YP0f/gCLq7Vjyj6AeFTBMbT43W9Us9G/Rxfv
b6jdAou+ozVvwo4GH6gSEPy1QOXVCMx2zhFPRHT//CbHzjUaupAg8sid7C9vA2mL4zWgHxFsAOM3
LhdaPaNlsgBMgyANFot1N8pP9OY0gQbNSk0rHSBEAcApg94d9S3pO61rbGwWcxCE579E9k935NoU
3uVWrAcY2Hz2yebrqHpmGJMonSeb42K2FPch2cD2c2eDHnxYshSYxtSzjQP0dfytpX8pxYKrJNYI
beFmghMGjopzO4UGw5ID0qjeVLdYmOBcY2s67rDdF8m0sgE+k/nGhJP/z38xVkPDkv+zdAwTULN7
jhl9mh3rYQPUnYWrfGSfmgw6RIvd8CcuaxTMS+sWwIdOkC8azqKGcVn+sfbi9KNn87LBnhv3ZASh
LskJWYYkYvqMm5t07+gYvrDZW+v9jv1HOWRvlo453gngHbADKada6FSHdxkOQDDXPR2Iq5AeFufE
yEHniNbeiNjl2mOPrxZMZ6TRGlrrYJ31svA5r78AgVeSVFbBpJ8cug7kN2KUYwNRPhqu4C2QmuNS
3ffRzpV8Nq2y5TB2/OuiV10M8A4zgDajhHc4nEfnxCEI3Kxey3VAmQcmfE5iljOBfO+qRIUb97u6
hDbkmeODYCX/RksnwZVeaJPM8KY51yr3tXQgJ4sa0aMtVpwPYYegrg1j0zQkWYgs2N1tpfWYNpo/
3RrridcGCWZTqsk4N8FEdte/Y65Epd+SxP/XRi5UCP7qtlB+lE8HGtMjVwqTcrkgbEj+3iMQR6Ns
B8bzCq4ayH4DGopM+Und2FxM1SiGhS3pMIsd0amLUyDeZ7AXFSQxgWxKo7oev/8fBthouempjkT9
9futjs64s/cUZTd4AcmFRasPMHot9TYO2ieOtEWmOUhKSs6uHjFyxJVvONmTu6wBR0eQ2eKFBESH
eFuMIws1icUto3QD5sX1BtxxQzVjB0VJ1tQgVyCvDKyoYZblTrB/1ZTyUDwqzEuvutZdBNu6oUCx
kFVObhV90eq3t/22NwM1N8lJ3ytn4Pudd+UxaKoGiST+V70kcTh9mYjT9hxvcRqoIhGpn/gebI8f
Q4BINQX5VSTrTYV3zuZL5XG/Lz+FjdV+EV26WRt6gKb15z4yj7QLrjmcaNeVpA2wlXFuD/TdSbc/
5W+5nVBQq7EFraGaxGPOmrNPCOJm7xETDL3Gga7EFmXIjwlmC0ftuccBAC5SmRHCrYIdIcEDp1Dh
hyRxwxKKk12qkwR/a3w2FTLlOxlaoA/S99sQCRxK3kdzqCSVAmqOrSaf/PP+P3l4S9mszZZBWn8t
475Pol9Eun/bH3MnJHRSZY+ngMY2nGMmtPkjiajibCcMQK+95+tYOoC5TDA6GU+tfIQ5zuwJvaMi
F15Nx8+KKkIYi2qmSup9ZMvql5lFpPSJZsxQLSPDUEqd3AYyMcMdlrx78/wup+ZE2VIxAfVqvylb
yXFRBk6CvBKhnZXT25MMe79AhCAsknYUIvtPyS092SeEk4THnxoC+I72hXViOI2AUG8irZY4tcbC
vjeQvQvD54i4VK/CinGWJCOLgBwP0y0n22On3FHTXBI3/vmTZP9p+bdmPViNDk7X3EedvmDioVCt
6DqD37vGd24lEml1LtXt7+kOSmyhODVyXJz7uiFmDBTL/SVXNjX89e+vau7W01a7pEC8gtMPKTBs
BqNmQkDJk1m/VPTHlrHSbnxS4N8d0ecc+uC+5dwZ2ALax7ZmyTTIpckYe5hk+MXLJQfIQEJNz0tk
M/nHO3FKB0sVN+u7zmX02m0AP2tajt9EAJGDsWh1+W/Sv1HGwqvJFQJV2L5lOuuV19x5v8YxqZ9e
PTef1E6Nu0bhhau6B1VRcrNJOcQdKBvX1T4YSsVpBDx5oNufcWNe9ZRnWHRDGHbb6nZuorOwhJv7
ye7PTEw+f4O0hzuSI+lc6tGO6Uh+0c6x+a0Y4VdKIvhdZE5xBER8XOIejIu0uTLyS37a2k+q6qqw
1GJns33B+q5Ty7XKqlk6kkQbnxuaY3xTnpZ/IAGj5aVwlG4HTO4YzdlSfHUkT1coQaZCFCEIZpwH
N3APk94m/do7ZjBxHsxeLnphrNrjJ3Gb2dCZk5FIaYvj4Tb4PSjAeAsfG7aDLdauWs/EZ5RsbVly
+Q7J9Ov8/C+y1tocjEMMsL4il+K3GHbASiInrAIf5MuK9MpfHxagJTL9G7X8+3QHLZjjmRLo3tVI
ETTqBekUGcJdv8sw/2NLHwSfRzHqL2ZRl/EabD6UUwOi8cMWDuURUaAX6SS17bO0/nBPC2lxsGqn
gowjxfC/ZPhF8LS92MNsRr2ftm7s0L/ylfCdqLm81N34RtPwuGFQrhrMrT+6NeixZVdDmqIfIkeT
TNSuJ6pbYIlVjodfJpWJOsalKbSdFINSzphv69SQgzbhnCJTtFPpFvBwxSSEGrZ5eKEI2XM2UjJZ
FLddJdwMq8bBrtReZcdSJUjcQ2nMCjwKuIrNcY6bfsjh61aUekX1qZ2AS/UcHuCdexLTZ+d9P3E9
ZtRCYiz2A4QnQVFkNv3Y3FRMPJ8xmSl6N3F+Z1cmNu9qOQFOIloWx8n1rRPYPeg9Iglml6tEfQ8j
7ei5KLNuwz7Ix0kLOjycpgYNRKU7MLVrnVXbMevAmg9Rj/bkTfsCBOJCt/LjOkOSBCHKvMZE/0ya
RsScaeG+wQrn/T43lvTMRC5IiNeTL1qwm0vkYxSOmn/aWk8YAxa3Y2QbDKWxYXPzYPKlCNjP9bxx
/vX8j+wcuGDBjbqm2dNLLJwWsgE/R9qq+K9BtugBewVbaxK8lJzFJOAQ5UksHrOi6uUB/kRnSZ7W
C6BZp+dEIzf/7SzbkIicKnaXfEoztFBGULl98E64HESH5WE8PR0/MJy/LyFlGEy5D23qbr1eMzjK
SGSyTTfyMYTR3NjPLRgEypA2/tXo6yFd+sgAn+23op83cNqcAJoSylau2xRVZHdJcj/WjJvyQ8cA
8ndcbMJ4bTrXtqYP/94pdLRaXJ1rH+Q9Bwt5geYc03BmEe8I4EMSVE7D2okiM8e0qofjiU5NBVHa
lNodB603sQvwdK4pp7EN+LSRX2O7HvIl2MCTAZdqx514i8UMhjopK/38W2PJ1u+7hMP3fCSyRGdy
wOy49+G8+6OYnWYSaFAbhPU80V9QrMyARBpcyusImKE3Lyhb9/PoCVkbFYtsc/konVZXu3dt9TgA
hC3nOhKZ+IzMUWTg+4BRhP2kQc0VrLbezh5RHrXub6Q5ixzS5KXpannn0nn3JDH2dJXGhcq8cz8c
NZpiB1AYBIJfXYAaWxF5Px34tfm77cF4nJVLzpQazpQkOqOPyluZLUV/u/u31G5qMf19UHM73l85
fflHZkssq/vHoPTUdGeOIkoe0Opt9WwPYp70TplAaBrU73l/1/hznV4oRCYCZZy+8DMTOgxleWeB
cfaCB4dyAzw0hhkCSJYeSjc+9ZQu7Uy9zs5GAJa6qPYPPVZxRm1kpicnTwIVT0N58Xy09oIFiPHO
eijM/zXaZoGOJgmT54aKmpzeT0VJ8Ks8znZfmzqE5DpSdTRAXY0uCS9quDfub1o0MPjjYsCo5E2m
L4fakgVSq0OXfHFdgpJQT16aKagucSClGa1sBWJemE/lYiMIijcYRtxUkdsWsvm8IglFSWlD1XPT
BZEBrQ83B4910HQluaT/sExpOrw83w55j8fb4sY3PzZuv2/NowpzyfFS9SrelvuiQHZP7Lvgjkb5
V/U4FlGqcCfSJ7ICAG1izR9ACZpYA+GYwszOzZqIfCty6r+uc1BfF460Ctjo7ovQfzkpem86lP5X
UCk/hH9KiCRJf0hKB6/JaEcqCkN2wt8XWt2fRYDhgImTHqjeBw8D1cc8crbwHePpFPz0pWaftFxr
L+266Q6Jz5ZYfJY+rSGCNATfCDOT3Yo0bHIaVdlWyHrGFsV3CIuOKCtIpuf4zRJBNQe4tCUqgHCf
tX4mGoOPUJ66OANr9Au/HRHdGNfNctf1BxhhyjoDzZCpT6izM7FsjKZ0/tqCvbtW2UfbBnR76gd+
lmP+7S6IQY6+Yy+kpQ3zKksiSwg3pqOreEd5nh7MH/KIzTIaRi2I2e/njWuc/MlnBPU7COIuQOev
l9nVZyho/RVg84jw36cvC0dl4gv/uWFZBVCmSYdaITkSKD5s+6k7hNzSWzfVAVDVLOQKVKo2i6lN
ijCcQuvQcjca6ytlKDvmLfHYycjzcHB0wLZyjE+RBldQsubahRPU+Bdmk2a2D31iqyFW94u/MOtE
M6TKNWTa2Y7C2f0kXLLfsUh9ubf37Mc5yfK5fqqTEFotqzF0ZU0tJZ36A8VA1Xin9UQ82rFt8fYK
tcKrDjVdhEFuMgH8hNAjcafewkI/HP45lod8lZ4KMlvTeC6t3F2Sweo0lbtWCEbjTBiAQlHRA/yC
VLoI4nSt2U6rCrX4lA4zWG/qKKGJPyJytSM2+5Mxmdp+AXJoLCLzEb4aFVb4HoesWE2TksbzfFx/
sVJr22s64d9mI8pL9TBQfJBtiRBMrzvZg+U+epeZwZn7JgRLU/2fAaE3ierGTZ105hl1tEenX2JV
B6GS8wxIm1NlEt5ProjIxB3IInlK5Bz7zsoccix1e/Lpl1LVBZlrmWxd2b08qW+SV5CdhbmvHVTz
Xyyl1SH30jbrbddelqiV3G+OZlKunI12ib7zPyyY0qZyWUuZ/MU6MPs6boLqbNtdmnV2J5hWIpZz
DNlRgrFa4dWAwTa3s7JlTOHOe4Zl9BYibolQnvc1IhfWW6StjFoamqnlhSXX6bs5e7NhT55CG7aL
qdbTtqIRPX9rJNOn38ZDzbX4AZZR13Sq+4q4tovdqWZfAmfH6xnzDtJQpBqeuNddDMBSp+Ska9NF
U7CkPh5x1oL0NpSLBOd8awkUgoES0oKUCJ1UVeAs+Mh2IcCJNsgsIGP4DDaTyKXbNsk8oS7+vaeN
vHHE+P1UacVry4LZike6VyRkLNt7NQ1duxnUOt4djpGeKfxcPAHhwUlxU7Jlyu+vmSq8zfWp+E33
nJuXKz03baXmrqUE9AvJ5Fn2HuPRhotLoLexKr+jCkggW+ASunB9RMt3/cem8H4WDpYFeeG4Vb/O
nki6Px8YX1oEPlcGxmgblcN2rqGdGeymbpLPirAhDpoFa12uPC8hCb4/4gr6pkv6x9GlHPF0Uovh
qY6IXAMD6XyF+K13o8leF+xtqDwCjLduKzbIn/qQQQVteVxLC8BhGW6UBwsyle3W9nJA4K2Dh2ml
WV0nD2jczB7EdFeJQKjVNEokLo0iH/wGXmvI7uX4LTIvRsaVSpJqMT+uFFk3JlAh8PnFs3q+DFm6
EsmiS2SyuB9sO0D3+pNwqTqjSKw1vxSYLrFXDL502XuAu0OxfnEbJZfcsz3vdoIvrulcMGn7GKxY
Mstp4yhOk+SIvT70IONq82bbjQececnr58rt8P3HUHFhY8xrR03pJjbkZy4A2nYxBURpRASGT6nY
25u17kuHtSPfEEG5Z6fix1YAiCMfBDIlWnFp1+1zJ+Kl5r+MIZAEefINW0y4O+gul9xKfotcMDkO
9K872o2CwHHcxdKnxh03CPD3hW7ytcwZw4xhcxnod2c4YcmOyTbOAvd+Gyfn4URqGMsU4y+9X8Sw
QLdpnx3y00N8YJ5KTel55s5OtiGNHpPJ2qxDB0f0lhtmOP+3hqf9yx/QrWfL0uOt2GU/OKBwdThG
8by0g98CHd/aYTRbUmEP732hnDO8O82DKfrlkAV4lBrzW3V0JOYO+3jB3z/x/wNy4u5hvWh0bBR4
jeFvWd5K3ENGGHpp7fCg83hYUPToPfvWPbV/7fXVSmpi0VosQR4EGngrKmRCpEnqKZAHX5INUxH1
pdrYZ+RjXEjXyJDKQR3HwL/1FuXHbBkht9zvhko1MJr8jQ3u0Ws2556wTvrVX+Mi/JDDHITMTcmb
VBQPRxoyS/AroeCwunyFbVuozrlr2eTjRWM8MxQ9IkA32KRENAyoWW1+Q4C7SJlPt+eKMS5DvbkU
wq47nehL0Axg1r6aRAlXrmsCjh9ofIrEWY669ifD1RJMEDtqZEFo2A/ecWxzU8tG9/ayoRcxsOcr
Qm8xmoa++Vwae33983shQ3dwqGbAocrHPrWtmUw0hZ5V9aiUPeKMgZ3G6u7aRAbE1ClYgb64J7nN
4sEr5MqRRqGY8+9IgsCo9KisvgNhsXCFP38PO1GjTGovDkvf2LfJb/qQl7xFDM9ZbTTNgR9n2CsN
8kBRMWpWm1BTCkiS2l/TLu96/uDShtQZznPULyZNOPUHxqmGLdgu8Og95c7qvSDe1h43HX3PlzwJ
9KmCBrYS0YLDDUYlQskdXarpNwB3TtwwFnn387TLjwOe4tmxoeV/cU06q5RKEoZ9+jYJBBRCjBcC
D17+m0tOXACca+48gBoB3FypWBAZ0BGaH1zxLkWmiIQsD+2HQSgTUSs8aSjtdVIlmCyuG2xTeveM
Rv+zMViUDad4Ly0wnB72hPIduvFci2yQDIv4YtpA5Lph3+3GDhStoGZHmO3n+gvjz8h2F3g3tPQr
suyGPf78PzjNy0gTsaoWNI1LQZ4W0lrVJCAelw9nXRkyZieJjbw6zpOKFeA/hkzIKz6dqEWV+hGo
CBIcGJxFwbw2KW/oMJRN1KqoIuwqMm1PGoAS+lRuWx1zrI3yyzD5jia6ocZbrx06CRSQc8RGsx7B
fdKvO3WLqt6twsFFoXfeMpoT2/M2vWcbM7DJsZDhZClbnhB0Ntx7BJYOWu79UqVyN91djL5qHtoH
+PngQ+lWyOVAOFE1+uwBP/A6V93+UrZhtdP1t2DPzmjey7PnLINus1C0Js2HVeUgtPut7Uni5ol6
AGnSy3FSfA20t3Eqe8aTa/aHd9lqBp4f87oT/aQIAVA++DsD0WlnFijUu6M5Mis0ZKlLdbbZUOi4
6Q8V/erVnZ7KbDxmbD4G5FhdmmV+7A8S6a/YYAOiP9+VDoDEspP+yKcUiJD2x/TUC2gfUuVeUpw3
CCNKAfgVeHJygebzch2gAYGRtUdWq7OrqqpdF8bV+OnE01oDaydtUKHRkqZ+vCsUyZSaaii+jX1W
2EfwtEGLWGggnud9HwXK1sKyEmPDYKyEJOtPIcK4bR2jdlMfYp3cTMAcLOPZCSw0qWqV4UAfXZAJ
tpng1W1gpQirC7szvPnqPCveT8qx854HCTgGcWyGbKfzw9ToiBK8koE3kccXeQ1lXZjv7E2CXGuN
uWKvfdc7kNnzUG7S25WDLT60CZ7Wd8p4B4yBL2z1znpUVeEnQqyrZNfxHGa4wSw7qFRdXDWldMax
N1I+4NyFkpFNAbR73C4e4iSMGb68J8HJ3clczNgTLfuuw2vUE7n1XBwbSXQqKugRlcUqKMItRQDX
z8cPDnyvqd7TNFMBqTYGuGI9mu2yEkhCr4vjzAAOBv8XoIg+IkEthQwF9D1sLRUXsZGkU/ff6/Dy
FXbCFPSclC3D11EcOdjwboP8ajx+0HkXIs+9ygcW1OsaII0pgn7mrfbpimGNeeduxPpPtjtaAU1k
jUu0iLcd+VPp65Gggj7po55JBZPYhngn5vtCELcOuMzbwUpkql0OZn75KtouzxJWDZnc54u5scr9
k0iwCQ0rpGSSQA8WawcbvneX6ksa3sLV8UHCtigurwM7ZbJh0W1q1M67oN0sR4CgQbi7Be3gf8cc
2QThyTdTIhmKCxICOjg6BDNnn/Ei1Y5/2aDZxMSL+jLDw25siiLnTzov8EjNJzAa17NrIBsqVS5M
DiCp2JL0XRrO0W+54vhuaByTpNZA1xwJeLdThakZHmdAAq3UD5Ub/rETQ9bwxnJ/RAdKfRGuVcOa
S8GuANoDOowMMLKksIstvxz1ZF9ua+a8A0aox5J8vJ6LX52a39JABAXVxrn/OpLMOsX1tawT0mrL
xDdAipvF7AJXh/SsBWG3rbYYT/G+5vpM5Ym1uK9aNkqmrQkGrdYPvv4JbF+2Js7GCLsVqO/2unIc
bdlm7OgC+S0JDWbrizGmNeb+l8tgfNW+GYGe8YtWLLgGK7XZdiB/ilWsgCtTWs+mJCzgAXiEaZls
dDS9Xk0vgeBknTzpaLCzQLyzZeR+vL8/CPHibF3m7XKCniooi9L2e6zVceQaIUYxqpLxbTq3BRD/
n8taPbNrkSvMz/7PdTsoOc0BlQEJNTB6Rc3mA0FMHmpAgJxRbmKePG2b9FhhDQjWBIpvxqB/9KA0
vRvMif0cRowJRX0knFKebYEiWl0iNEkv3sveauZR+K0Nhe9bdS0aYiKJq1+pt9ea2qcoWZuev1YZ
I1KRP57v0iug98Jb0IAghlEIrc059Kq38R3wYw4GdeuNtMi3TMiZ5zYqmjEb/XEN8lViVNwipGJi
U02bfj2LzMRMx8lggdfSpJ2lk0eCHH1esfKcpqQYwCEPvYZg4yNZoE6uDl5SUGxGApFcoT8VJFsw
6STUDU9BTLuB8F19V2In4xt/x5kyt1dnBeHK8CjLD2uSFR9R1Z5SWU6qe1Ivq8KtMS7sVxxvbv7g
ucJgbUQSxmt6AhDUrLvzZQkzMe+LSRwI6/JV151esp7wuB+mKVPOWo0AyBy3SXVcOnFiY1ZcCK9y
eJ16IQk1BbmKaxv5KMep65zZMIxkbKo06ilaWUqHwQqlKCIHdHGjK5mjP/LpVd70U5u360VIPaVS
bWM2u2tojzZVlvWJGdF69524CYiedY9nj4VWyYNaHaTe54nOwB+Rp0Hsxe0q2q72dLbH7iW1LUCR
P7YBo0nqy8/Ij9aBpiGV18L2l64pAEKfK+FLOGXWYsankPHiKk8dOrRJBo/NpEGQFkN8xiQDfqEC
n5sye/O7Ex7jjWZuERq5a/K+oaZa1CM99BNZnCogFOwjxaILSdVYY3KrT6VJAcfVfTs60CXU7KLu
1DVjIXzxGocMKniOuZTPgnEq+lgwmVRxLAOp7yoxttINF4hFyCYuU2yWvW6o6vXysJ3ffyec6R1Q
CZhXCFd/4d6v+JoL9sx9Y4vnalA0sVvwx+z/2pCfBqk/8MEscNGIIAwH//ojSQHUsIQgRh6YKiCJ
YvsdLpwJwLL8fYpzWCJ6/nSFEJKtGbTWDmzWIkLSv9lNcYPGNrvKh22tzzeiQA/rJOyVyjkXtwZX
YlVKVW+OqPoZtrbA1/TJ2FosYgT6cH6D5Swoh6oGbfPWiJezlWHpIcpv0WuSIHGEMUAxs3iHRt3W
6orFUxED1jXR7jE9ytVvnQQGOT5ekZSr6j/NyFY2EBjBVeRvkZwhIqgmBF8MUCHZpEVAjw4nOAZ7
iFVt8B1Aq2JJ/SFTbOjOpFgxAE2UEe125tVbKCFax6mMfQL+hNG9vNMt18WIYlR0nVqdJDX/Xob5
XwnmeiDhuXcVrBEH4zdw/3wt0HMcKLfSMMaQtFfSuK4UStyzxZdfwjsXcWX74oUKUB+CA2XPgtLz
nmbN4En9G7cdbZw6RKWH7nIxMJtUAq/7DIvUD0XcFB9+sjxeaDb0DFR+X19pycjwiWbEgAo4frUp
YvWWGNPxWLC77o7Y9NpZal9lIfTNfK8+vdPFUDA6hn/dYz1nqQu1ppA9bwcFGdz7lSHNm/tH9fQJ
UHMb7l5ijAp0qgh/lzZcuZ3MmqNR80Va+LtJdWaFpkwyhhinKY69TSGstAQ6puR5B1CaFMcTOfDz
q31M7b9S/8Zd8kMvfPEClggMo9/Qx5nG0cN+ns+pJCIu7kstlfSAvmRey160VCxGBsTpGfbG2GJz
JVRGkQcXe5wwh/nohyrgB8Mm72dsig7qnCph2q/Zv/GNkOsrQJmqG2L1lhmAPgE2nkZ6WV5hweb8
HRw1dDfjFycqsxhz6FkTHTuxrdH/bvIox2R1xzjpFoQb/fJTbkCvLyaql9MxouGM6ZrgC2v7rzwW
FcYANrBXrwIb8xOoR62NQ+RsIh/ZIBE9HHwDdDbn3dnhs0Tvum/cuK4/asEQC4ZpQauBBuKV9lLC
SjAw/f6/NQNoelfX1/6dyDR2InvTRkFWfPk7sRPtkHu/T79DGsBdz/lAwH4BBU/xn0/1y6SVZtng
+wUMuNzfib0CJ+6xaR+FkJa3GOyhRXYTYzJzNQ3wAiTqBnlu1m2Jlaib+eLYgyZjkhtx3zJFdWIZ
nQ6bPxtBZF59gXm3Uj+7jwydv9N+GJLH6vWNFoqRd2dyBuPaZNP8RXY+hX5R+DX4CuRIHrRsW6rA
xUVYms6InO//SaPqZ133JYaA7FWZxWuih/8/lWKTSb09mdpFVFeToYh6UI7DOmizt8hxAErTXbIP
v+oZ4CnhiGqX2FJG5C6tpJaZPEIyvYgUDXh9kUiTXN5opYqzZtnS8ugmO7ltAPT1ZI2dPo1LDn4n
RhIsISGs4WgbA5XnN+isc7X87x1TwgqPX9M93qpxH5YhVZSGpB2mt24kpAoKuCN3E5h2fo1DOrRA
NwnQySkHYdCyzHHupZoIgnum+0GWTaOnSf+KeMqJlDCGsHWF0CwQSPusi7XPLFQR9HWtu3uNIQ7t
8dBNiiK7PIEe106zSjCpS06AFH4Y6LBCnqsxZmJrWK74c38DY49COxdTmlb2L9TF/Cr3e0MygYRq
M64VurLkqobRPfUnSGBWKAYtW342ttmtDAotRbnU77EnNPhQTlx2ZYxdlBPLY2SoVx+CvjzX6YBo
oA1JdREiUh4bgr63b0UymheDN4eatY2ijhxyctY5kZuCmuv7uMbHNjQhFRQCqy9fmE3ekkkkFd5N
iE4UUAIivKtQXMfEI72YcOZbXjNyrjsptMl7emtc/QOFrlJl4GbrBqBwHjCe9/zieSlAfu7XnRT9
sCwplVzgg0/KmgUKENxRzy1flZ8pJGVl7E3HsTyX61kkzG3r9ShoCeHHOZKTcoNzKoaRBHTh+NWL
tlp8sKvEI02xQeTi0VWLSvlF1v54v8qsh/q6+V+Vw+fl9CzMtaJxW6bzBQ4TSvRA/oSQ2RMN9eV/
mV93ErBC3mwVyarIA531w5t4xZWrVs7P6f4dkIrcope4ItpEBC9wSyebzBKVbNyHeMXDgnxHK+Uf
09zjCsrd+2ULvgUYAo5LbnKMMg4hY+D6jB5rbdsTHT6W6h8QQL10NVM4ZoczkEjuGVLOWefFzuvs
AzoStR4Rg6vGC5yB7A44Eh7PjeMORxa50SfDnz+YUwAK46BZriBFYUPjmJU7XBEQmoAg0HaA/Oo2
uKHIK0e0XJQ6w3bEblIsmKQZrdtAu5ldkaUpgU5ovk6WSJrqsBHXm0nD2iYyyzCoXguX09QhFfAF
uT9h8FwSfL4IwkTfukCg0kggDxGUUwItSKzKV28YRwEIW8sJT3TBRBroTaCy0jJ8ECMDQmJXrOmC
dyQYJm8N9r2nXe0o6fzdL5Jp3SlN2+kj42xQiDt1ceY4ETMchF/6uq4jseIFHFnFlVw9mV7IENRw
vc3qJnVAC+focAo1bh7QUoBscx6K1QwxRjILOs3V0UFtmpFtXXPMYCyA3fgyPnVQCO3xic5eDOQC
fkZknGijf+KCVvyn8lnDHpRw9yiBRQ5eYtqsUoIF6OUEsIRY9uYL/yYAzdynhm3AtLMEIrpWsUV8
dh+gcMwTPBVcEXwf4t/wM+FtMOX3BdSUhFiMYzlyrcth55VOMn4GyjlLB7Fk55XL0XwgNsKo3Wnm
58nWBNEIfK+XdDRrJbXdgTAZFy2bgqZ4zcGdSnDy0xbs8C3Yfq25Cz/DqqazlskxWg7sdF5Unhc+
cIvo6GnRrqAEf4t37br4Tj1p3o1biY2s0gbubwjaXaj4wAt98Db7R/kyPlifxXTnbqsT5I6R80qQ
SRDnFXxvDKYElRK2SlcpJ3guaaKVesn2inwSMeSxk8hFDp+tSMmy0avUVZoghSkiYqMgGamLfSOZ
aQ03D0iurFnZNTYugLjnBJjYPuuPgr/UADoCnUeQzQMN7gE1NSNAENVRF1hoYKYkLoNGWoaeTqE8
VeyAulxop0YfqCTQXkHDc2+zrDT72HPjurzFA5sxpHVJ9CclF9PlHiYyp3TQG8w69yCibOgAqJ5+
kjMPPVznYLLek6Q3dhnnSlfsx925yCa9hPD0QAoTw1t3ScH0OAqxehjqzmoyRAjBSH1Ej0ibfscC
uEEnxt/+RjIo3evAc5UWHay+GfEQUdffhoPlRADT4zfG2IZD6z5+2qePEKvAx7F/ALmzsmBPX8WT
SHo1AqF5Vy97Z5oTf+nAOkpEaIlZ3XGMc4Ac9IcPE6G1hch67/r2dqTLN3cVQP74OH+4xBmoFngE
vTeuZezWNoSrz15aDwDNtmHyu67QfH5TX6tDPj1XS/W1VG0vm4z+MyNNIqXgBAvX0aVo1UmYRBuQ
bF2MQup/eKQAH7R7nSlpBHBver/Iyw35hybnDEo8otA0GEzvD1hZhfh6JHwCcKsGz3BnhL008fn8
7OeAZmPxDekwE8D1fKv/gpJ+wOI3vjQmf38mIt+85mZswwia7A4Q/zI7r6cfvliOP2s7jBZz7rBk
Jm9SzrVnsChJ2cpFSoubjfwCPiWYv679ONTUeHMF/PJCtxf438DzFKpLPQqFxCeb34Z1nqs5I7+/
pGMgqzdZjcp2V76dqXpHGuvHptr4AYqECWSMM3Ni9BDQwFkK6tUXD68CAj9FuXK5V0dEcXP2ydCZ
NhQJu/VBFBxqoGuzhrctrrhk3UmNBZrb8WNVb9IVu98bACG/2WqYu0FOUzdh7WtULGt5TtgKo7V0
de5N9bVkXeg/HiyIhyes2c3YJQqdB1RrvL45RpIbb6kT20UUu4s9j4L3FFF4xRvceOJGC5+XvzSv
7hT4L1XHIKCNh29sPzXikMInkVqPF4vMV9NLyemH0WI5/IJUSI4BiSoBi4q8mavZxHhuXW1sUiqH
2tmvqDjn27JCOVa2LTm1T5ui250WLTKxOt3TNCvIhF1zKEU3T60BncY2mr9v3cGAazRkSQI3+85L
PMc7XziYf5CJgOlhjZiAII8XQgamDJzsF1NOS4GCkNj0lcVSSgzzBfaSA3DbCxwXXqOzX3XTjFsK
QzbXjiRZL10syTgIQ0nrvc5iHu/Q4wLYz0qTkavuA1E9tlaiTuRUb1bKB//9pXprgcOOeai2tJrQ
3WKSpYQOsshNE28LMigYcgnD4J1i06CU2IRGBbFQyBpqpQxX1RtC2BONm2V0gT+2jDqD+eLVOgpS
xJExgjDaDfFbJoV7NGEe7XOUz2Rt1xW+0x89kcCWhiWsR29CN1Jm8ZJrU63SEejjZ6LH8BISU2bJ
1GFuxbGfcif+8F3iAGSoL7ESBYxYVhKvade5u4VbYN5BWDdDmNhoBNXcaqti9xTcdQnj7lBTKH3h
NWfqbVdqAtU/v2LarsGDnJ14kSeq0NF6cvfVXn2Pz6O0pRA9l/u4r4rWwXZz03qrNDOc9j6XwBZw
5zbU7ScVaDM1ZyGb5XzF/fjjAfr4zszG2UDTXNmiua3cNLR2dwTCfEW+kktje7DJG5caYFSIIkxg
PwmzEwApEyc9L7+z2DArf0N/m3ifk48uh/0HyNSilDQKmvybHSeSVGQ8+xRMnZ3VGS1N0njhzdNZ
pAg+cZKquXkK0JqbTpIljCq1JTYwlbCeGiy7K2vketg1X+FPj0PlwE9Q8pgOXSyPxB8EoxARe2O7
qBdJdKNb+dOdP+7uqWk24gnRz0VjGG5CGi+zF+1jbDnzO3KwQFwsN1e6r3u7K0OKA4pu+NE7RxOK
51nA7rXJzS32bg15B5VyfzPIoZt5UI1oYrKlcCc69vCrgOMPyuePfXWZw25YyovhJV+5ogAElZcC
9xRrKSbq8Y0Y5J9u7GBJhw/4fqXQQo1M5ehKkxg7z5pHj+IHijB1hXINMhbiNie/w6+hmrXAy+bW
BeDlj8ix3x3Sx/bPl3vD1Kjfr1Z2P2jbHVgCFay/U/ZZTkaAjQY2tme5g81NL3Y6fDQ6kd1LjYXB
qtpKBDUnjsUc4tuFOK0Z3XTsMXzBXCsZBp5fVdVV5C22a1pc/GUjWBQ7+E+cfhKTRHY5Uqbp4BIF
FQhe91+25uobPkB6UnSYp4+z/SzPpeoOHhtv4MQSpx9yYFXROJ18U7Xsc1loMipfGYQtmU8NBq+F
fVZQQrbjbo8UsWDP81zvWnrddwa+1TwcMJWMCZGQv/CQbsaL8ZpWSVo18glRqZPyOsxpInyGV+wX
cSoIozY7lAc1ULR7l1JjaCet3tx1+BsYeD+3KxZlQWqAcgpkbHN3TMQKMzPCMLw7ZH5rRIxwTx8j
yEqzgDk0cLtIw6ZZeEXbXIsjILU8NaeeaTwbOVQLEzHueUjn8aYUg3+fCnfsV5q6TTuuzu0vu5hB
PZWjrYfynKAV0++4rxS+VKmmyEP0rMUDByubY8slCBE3fXmOU9nZ/c2GdVELJNGjGjRsW2VEEDwb
4/SDDcOy07B4pLAd3q6JaI4rIu2UnRApsxWr2gNmdnmKTj71cyse7j5U1eCQe1iaU/oKElIecU9d
RfmFy7/uWLByQw9VpV3tXl2rn3V/ISauHJlXxXWw8boWWMK5lE3+p7n+u9sCJZRp7iS3sMa2fiQY
uB+I7ruMTWWrFZwAdud1fI5s5bXXGVvOeVGUe749plYEo57C7SpPDsaqStnDCmB6hQbSGrGaJDq6
NofqqVRGNetFf51+FB3HpISEL/+Z7OrEO5dBIZPVZI3VbVobTdYTvgVwC6H1ZCNJ66JzgXkrQvoz
EFQoVpXRWRetHIZD7z0ayuA7Bz7zwPfFhYfCNN/wCVZQLJUnW8QKvuE59kpsZovqsmzhrERa0Afg
MRXdTfXDXIgS0BuI2ja0E+90oQhiMPWRi5dOG8plEtYC1ezEkjEvIZCpIq5UMr4N7sJLvSjZI8Ra
xsFPX5IJztAD6jxj/13y82pK7znrIbQ0riqPPFWs7I8YKVaAbNlb8awLJyBVIMbHhAFHfgV40wtF
DICt+5ehccAeDVClI6rDnLATgV1eOxDNHQaT5d3M7KUiMH5hq5bx4AKVM6O+4KfR/p1kBSLyXYQ2
XbI/JTsJtiQQgYjI6LnT4ingMTNlToip++cxWFKy48nweLMkxqyJBo9IwTvUeb/xYnYIZmpWqRi4
GRGTiTrtr7LYylSIRJpvApCns/iuQh8hdv2PgABDMeoQZI89FjRbeVa1MaFNCO81VVnlTizzrRZt
jHnkdoOgb6Ba0qOi6dmZeqzZKOeotoFHtX5RP3PEUa9ah2M5eYChuvCOkLOoXvU8YCzG3NTKp90A
zURXXLntU09P+xYqIIFYSGJnOIl3YDzjmhWU5k/anThipCFK0OJwyuTe1qT9RaQ4wPhjoeeXxJbq
/z48jJ/8aWKPlPS6u/Ax1M3guokrklm8C/UMaDROJQMlozRRIzNXhZrcY9a92TzSK2K33ieFMD5H
lEnV/3C3J1bVmzFF44ol3BDQNwmploYkGbggSXj/YiXfl8PU1G6gJOpu72GsBuK2sgFaYbSFXcpc
TfjPfPJYfYUiLLmBDwyNIU8iRG7IK0BQviZc4vmZpl00vzOg3GvW+VdR8JTTTi1F96B2+H/4YL5e
JweOT12YHZOKTfIhkaoOA8KYpP52bAVqtWbGYCVL3rihnAJv5R+euoajzgNyx13BUU2kFudaypNc
SBo5YOBNxLRx2i1Is2pSw6UIUdCYdH/2gp1ag4M2YojpU6o0tp++hvKn71oFrbi71E5khVedLhe9
Z3vWomAyyz2gmficU9zJh1ncTnMNIcSvLR10/X5Kpr93dVFvdh2x/h/vsnqKOCGUFbqUvuFa/EJd
n39LIbS6T0CONs4vqoxzw8xrfbS3zBYHFcdKFBtkYQ6MMrWkPOP0DEptllOoUoZ8LmIePmkMD9xp
ZvP/48owU42cLojwBAJBwqXfLWe7xDic6qfMvA3Glc8I20ZhYSoV0PxeSg3B98iLrES2Ke8edSCM
5Fj1hMDqM1lFLie+ohRMHifaLjlmEGIHYNzNQws06ZlqI2LfzPjCyqAJVZm+8RgppHJDbnG+2c0v
3J4UwuAcbqiQK+/tDDGlhZpcmkAvoz2ghOC3vEuyZryv0ttUOIJma8I85eUcrIfUWMu4hHZO5MhK
5Z7lTIDuh+Ty1jrLHmCjm+2UZRpIV8wi/5t8TOvjmwZHDUpY4sp6oZZkcXs9T8Oov4LWYoWGXFsN
4HG7lieDtUIx12I38stWEVlA3d8J8hQHoC+ZxjrjXTz1SziI7Xm1AsaN9iN2xpP0NvDbFQXmpiTA
p03klLNH4KwZKOeqW0n2lLbRGrz2G6WbLzdIadGE3Jck1mcOsnEcrKWd7Us/PpJTaadLxUlJnYqb
zHqqXBA3Yln3aeZ20gnItJTNrF0XkDZDph77rj0sBaH6x5liU1GhYyD+V1xm6X/E6dT5i0z/SL1U
B36NFP17ghfkOv4vW3W+CIWMZNwoSkRVJjsjg2PYf3RtcwCWX9n2tbw0RzA7wmSzHwXSVJNXVWhL
0pn0ga2TblxY/g4So6KlkYeYcMZrKQOEfVhB9dWq4cXrIm9W+8LtTHnfvkddIanV1lLpSc3eu76G
/SAmPpohp86Ijim0l4ybi7YP8hkEwilj8cA0QFWapsplHsd016/+r/cdZzoXpWAq0/WgAMrzrlPj
iWmKglNo+bQ+Dg4HYjlt0JvTD5PApCM0qFv4PyJA3XPQ928h3/uA4mVNjfVF0UApIo4yU6K3rg5D
OFfgSNRPDhZCCDuXcrgO8fKwMQQzOVX6qRBnHHDWn/TRruxO6VbD50QkbGvrblSGR9QgBucC3Q94
pY61NZrSta1OVTW/qsMOO+dTInBE4z0EJN0HaVTJVW6o23RMf6dST5Fy9ic16XQu4waLPeISdKYL
4txuuUsJEBrcWkMp9U9xPAF7u4qaJUtitlc+Z2FHLkQBCOjFSE8ytCVhMdMErwIHWxx7+aOsRD4n
qY39G6e3xhWwUxd/S/Az8bbazqy8mu9Emg+aqQit9ONLI0sLAqtpJhusFAXUISJrK42UB8QDwMPY
JiliANYcZWlzkvDwSSF+MQ59n1QBBoQrbqN2TIU2jLIDEkp+iGemhqHqSioWtn/QN3p6ivuu16Xf
tUFyUi0TVUrlmwUa4FnvON32RCKkR3+JY63F8BfAJLBLBCBpSfF6xR8hGbsaLl9pDGDrxRD/7GEy
nqFBk0Qc8BuGwk5vUGcSApBVHclHcW/y4GlJJ4iJSxnXpwnbCtp6wNZxSQfADdXE29j8ni2EeV0B
8YHesyZyrWHF/LSPbhnOY2tBd6ywmDOL0yhYinsM0HGop5nO5sDs+reylsebb+7sDzzTHSa5Dg9V
232l790nuTN+xLqm6Y8zVuVCWhAWg/6WI5uzOh1lvRKu1WZB+wivScLCfryfnkZ6g1a0pXSl1y4U
2IoeRdwPtH5bNrsuNdJpsq8z2WZaviEdDQesg2RA81fRV7T3tGqLMlhZpxNEAQ53BG2HVuxpNPhO
Jju7hFvTZ+dzn51LMoqemO0oGXrzAUrJPWk5wa3x1IJpDah/bBb/nFPuWmiOLGSCJnGRuv7YAVMJ
wm8Fvf58IpDJHkMJV00jBVlbCKYWePasioUvPTUa+rQifX3DS3Y6ETwX338mZtJTeY9qUiOpjTXT
yxwIFO/oN3/Jj21ibOu/CTa2zx+Q2T5++nLRo1HVUSPt3VcESYWnWK+jj1mq9JRa8xYgwWsYERAV
fmACFul+0STxjdglHV3rVvsZQ+LR1G0mXd0lo/TOAdUnI6yRPmm4K2eZSlAtHAQiciSVFRWDDs80
QrTb5gbrhPcnb0SP+5pJyZ2xYtrk6x3+A/1aiEzpebaEbXUbT/UmI/ULi+O/MddYIcxjLohV+OjJ
HUu2RHQ6MQAgjIGnaZOcRqDOEuTvbM9slLygmfxDwv2GwMBPqq6USYgLL181ly3qh5swb/Q2bkEj
Lnmm4oyf/2edXBWWsUQq5SlFBz+FggSWsk7CRJ+n8sJjSEdiEsw5K1zulOa3/E5k8KinQ8Jo72fF
SwL0+o1rt/U/KYbc4ap4cwpEmM3v8FRHw5mTmHJN0k0EAY+yZNohCPVdFjbznaO/ZMv+8612Mk9Y
T4WGj0gPbRE1oiyrg73BmGyRBFr/0ByXsyXQJ97hjj8bdBf2zwlL7S5bvbHkFpHdGVHz+3P6tgec
CuYD01Uc4bUEZEMCTT8QJrLvHonSBMWghqYaPzK3FpTTJo3c2LtFw8shx+xFHTViRuQLhwyAJO+P
m+H3rjryAztXOP59Y0eAH5VpK5Dls+x95gPr1fbL101ZnMUrL3H13gsDk7G8IRdPTQNLkJV9ALJ0
vETYpxrmRxzrjQJB1AeCjt7HwB4FMkYV9MkQqBgAYYvZG22iyWz9PxsbMVciBuI1ODrgx7y0Nan7
tb39QEUUvbXVSeQXKuHvq466j9eG/HpiwZ9PMZQeAUxm6rZT9XylcaH/Tr2PiWuMHv+z/aa6fxRY
s1wHzbqK0S3ybnkzMuQXgHd8QYpLYSJnXf1rlH9Fim7zuEQA6vgccwwJAi0yxHhImwOXA9BNGNp+
tvxdcILjG5tOO6HXalUe5DPYog7bSXGy87k/i1taNdJFaXdlnnfXquk2/2Ibe5gGvcxKw5kpcFyD
K6d8ynzibtUiM6KBP1etoM8tc+zQ9tLSua6x/5ceOQJBaUnkfboHVvrUYn5VtNBDULmeCaSMXe7e
b4XTJU0tcClDDqzezK8W9GdwbACby2ZZvT7b+u/3U3ypl1uvpXal5QgHpDjOOjAvo6OLigYlkG1Z
huoGLDl9YXFBTygVyw43HP05CpktDRZdwuAnVi5gH5q3OrnWHhYOz3SxD+C3P2SP6Wg+WLLC6AAI
RniSoCjlNZuhQUpbn0Uf6Gk75gxZwTQEPMfGJ/GQghdXVeKhocNVATbga7fU14/lv2zD2dRp5H9p
Oyw33Pzvl6etHPrqqvbY2gg+jdNJB7WAhCRLSVgovvCW2ujtkC6c8tCW7x4Tz2n7nfKTSRdNafSE
UmUMLx00OVd6nMMpdEKpEAtX6EYjZfrFbKkOIoCWTV2Jak8a5HagPWUtRPVd1Oiei02PoIfkmQG/
a07RPXjdaLQPOhl6irl5wwqO1PAu+URfZk4B9JrpQGlKroQQ2hqZHI3/HLGENA0rbctR50nN0d1+
+5RfryWK7d5YrewUQvZYKefkv4jJGRx37rNsWTHtKhR5bWB1RGGLfm1qOZkKg6DERQ6CxWkYuAIk
v09JHVjlj2jdt9Vg/a4zM9NdGfJ92Cn9QazNwZzUmtNcCBqGBMcGSdgHv2pWTg0SNxjBi+W9K8oz
O0qMDjcAMtCS3qLhvkgf9t6e60iLIUrcxbz9KDtaSiFp1MFHrAuEmwSXpdMAWY4m8MaEPJv5Fjra
Uo/NL9rQiQHV6rdJMAmey2LBB15QoLbulr1BI/JW/epKew4VyA/0Q5aTc4t39g/DcoRrS9sQ+pVo
99+P0kyoUR7RKEgZiqAoRXv3lvqn4d1jUyESKdLHJg0CGYqQ5LtaBgB7sY2fy2GnSl0gukPZMyXw
FPflHfGc0xvifM5JJvLw6yYkmTm8qEF9TPjNT7NvXsCCoRSKi0iRrkzseGAQI3wU8ypwKO6GJS+w
PBdv5XM95cupYXT38T/VjUL7afXcvH81vmgqiaoa+yAP1aORVoPY8+J+bwm0O+adYGWNlGgqkqFH
3FdKPTurYo2oF2VooVkAGdUR6mrFIM1/m4Zg5d6ka4moLn1iu43FbBpeCZSTMMPQWNwzy5foqksq
szzc22Oh66E1UAsmAorYptLPbh0MGP/phP8vAN5Hrok+1+jh6kCMFP3zOhlzE7iPYQZczPjtZ+Vx
vj39jx9sO15SGhMLclEMjOYIARTUQHj+KgYQ4MCTa0jIcXL6/5HYPZrNtHODlwqP113a4e0AMk2B
fjyz1BJMPRTUAr/POJVL/JSaGEENGDg15mjscuC9xfk19MDoA6cLvCAimwBkEpZvZbzunhQ5/Ray
iBXGvFBxbYyAUrJy/Lyu5AUYfQein3EuWpm5U+ZCAdtQjAKoJfl9E2mlW/6FSH27aiiivz6zEmcH
qwfxvYaaUEOmQJQifUKeWPm5d4zrSdS/VU4oCt3tNMDENC7+grkhcreBBGNq9yo0VUIKytD9h90k
xVfZbRiMyJ/9LNGSWjWiN8MvFfmLoGwlhZvRTpxajWK1WD3tU08FTEEPl86nFHE0Kfs3E44eVEl4
c8Wu8Ji7mcX6YZCEx+fAFKAS2gALC9zN+2ZnFfRG5y51MnOd5q1Xx6aXIyaOVUnNPXiXlX4n9OIG
BqVKcBS4edqf+jIIOFraGm9eVKhm1MmtO42qgF/mTnSfxxs/RNlNx2aBCIwHvCfW1Nxv1mAB8vYq
5hFzK6lvnz4BBKF9oypWPE9EZtuUwXZnfhFklqoy7X7b8r0OEzL34ah++xFQKJXNGkiHwhNwNWHz
QV3WFUOH1uUsJRxh+wPHAvntThUK6DnYFul2v7rl7MRL0YlXomMfXzg6mqnGIcq0T4eH8RJ1VBqK
JAtT9wuE4Vkl16jjS1Lcpd833wHnRgFnJBQPc8sD9gM5lnPbLOqTBl80OcqYjEGdonkHFlhg31YY
kjHUEfy8RcgZotoBBHIwoSuf6xyYEkcbp65bjRdhnDC+UkBuyw3R7DPF69q4B3glk1bS6YoI9aMc
Jal6cvjLOYXIl2jz+3kBg5CjQSDRft8O4QCfDnC745S2fKK3uoakfUDvcxN/ctbud/3DGCDnuao5
y+G9BpntX+tC2U7CTuQeFYXJOzx/+cLT8jh94UiFSJ+V8CdvIYI5S2KMxbZEOEYEK8xicTDdg/UE
gy8j5ovGAvMuGToxMMm50RH5jUPDkxfF6OEowx2B2Xj5eHbBwCz0b9QBmE6YH5ivsZWXyoIHd9n7
qov1u2dvSkGLQVSoHDCXRC6YJhhjW1jyMN9goIQdQ8omugLlfxRWn6SMmYC3Yw63IjdbqGRHCC0z
ekZC70Bi2xRL/L2iF07s6q9847FHK5+yoaDkOV+9AvGU+elPDaoNf+7gUSX6C31PlKRjQSZYDtGz
8zr5wlc5ynqM/9RHNqWQ3Jkgeyn3KUOGbEMAglbBcwnCOvZT8HI7eOT+YZPsek3ymOoBIx9Mle61
Z6/NaSaoTKAr610nc0aeOCG34ilDc1uwrJZhVABjvUwp9n+tXco8lf51SdSebb9IrrrqoEReUYGO
lMMxKGWbWAhRvtjxPdHFENx0YWyumRIMawFOTfJlE023NevM4F0+43ZEliYp1lAjOnTRkn1siHFa
ekl9JkUhaM2GsTl5OUqKQqzadUyjOoPo0hULicrGgQfk25v+B+C12Qlc7DLcPnjG18oI0P+N4CfR
FcB+2RNRdQ/VCSTxwlXMuR1ZyT/S5dD/LLXy+v4bXla97sCyfJD+065kkNZ2xiTFRMiYqpvUEcY8
yTRdLWA6cnCk/cSpjL6TAFo1flI0xG/oE/5Le95y57oboLrzi+AvJZIA1HMijp7KHIGUcYPW7UKF
+NUJPld/1sc4sQ7itlFX3m9WOkLlh+7CcYuULqPuOPonffhiom5L+tKSxd2L7qpvStktv+TPPqae
yvs7cZvmPwzDOH/6DexgQ4X8HQ7hbm5kD6KPIYbFQHwiLKlDCj1W56KMwyZJ+/t8K3sEKuK6a9zn
A0OObj+/l6hXtJxmFpyGp6coUme4v1s0Af/mXawFcLuXEoBI7Tx2lhkFlgWYyct4pRsrwK3+iyUV
8AYQRNstPbaSVBNWBYI3r0s6dOYNXk38jsLJnZumyB6r5iceSuE4voN286qyF0CI32CXicFHAq0i
7x+cjh0b0mnkGLEiDnDUEPiGncMSWqJJLs2vB3MQE/Yipg64Od4WkD0RrVwYxhaohlxmXiK04SH9
MIILTFavSl4Z2KPEv8liLYPdJ901mcEjBuWWgn0+afrfpjDGN1mDDFGkalgOS/5kEK5ZEywV5O3q
/TtMDmdS1pFA9dV82ZpMoX1ybW6GByN+tlJScYXGrVUq/dnStUlnzwrwFZYKiBNcGcM+OngCE1MS
LNwvGItuesIqb47Z/B6xsdehq10rVSrrKyzYTkDD5z8AIAE6i2jwSUGkvkGyJ0/hRSGHd5kJwQSK
OPgWNqPEsnvo7zLVCHdhsVtsB8haMrF56ffV9TtBGMXzR0/PwZLiVBy4aJcVHQebLXYBW0SZZOZb
O1jnyYJueFenpPbzRKOiWRtEFnDn9LdFzbByTiEO7c7D6fkbxCQml6SYEWUahmEwCwhtR/P8dp8/
LUNpCE3Erh5i+XEeFWX47DDJkTA56hPQvTQGPhxpvEC9l1pIK4Fq0pfUtNRYjg7X+AsDvoK+buUe
D6q0qEDr0/VKQZVSR7ecC5mL8FCB2g2dmF2WdV67pGDQoyQEuq/FPraABBGx7yYfCB7aw7JUhC0I
EDVdNk8GV3ni03mSy8p/EQI+NEsVIGmEmdrfp+0mn+A5Coww/SLCK0237EwLMP8h0ek2lUDscmaf
3NbyjOpsEgyG27yuiLB82ikFPFW/C8Uiacug2/YQFKFdQjwgrpydKNfL6w36pYAdj4kBqpfYaIks
4kJMAEFbY8v2daRuxXvXNXZ2oPl+1tVj5ihBFR0ZA5bvQdyP3+i5eVim+vOmONRbGZ0a7glRUcrZ
00b8V7vRG1YdFGudM3j5SGeVCDv92Lixp7SEGOdG66N7CTX1pNMbHUxNtmJgTVtTxg+IDeje1YH0
pDxeWjIS34ywVqSLORA9mvsWugJR+t+CRCsw7kQujUcHBv+P64oFrn5Ibg27FRqYuucPggmADIg+
roGiW8hAf1saxlRjJF+Qida4rsth9QppWUwdUfWyym8xIb8ZhVQPJlPENfRzFt4jjhHv1hGTl5Q6
NMF55m15ZiyeM+4GhJOhetwtICVTamwHM1F90eCbiuxyuSYX5VjCC9fkDJ0+DljgguuKiChwHHBa
4hIOdYIxnCB8RUsTUYdCN9QvNYdd1GPo3MtK+L4vxjFiPQ1ImirtwmQyjt3TKbm98PuuoeDQqlHk
/3nA7e31mZZAtOuZmnAFODqofq0AkyjTAUToVPSc3igawjSev05V8y+8jMgybwK0dtqeGTrHdOYx
cgcSjNVqVS95Ui90MxnNYR2ydMySTITXW4osb7kqgytmr3E12FYJliUxnbxrIjGa67Qac9qV4ItF
foiMmYYuGOdBN7B1wHbDpOQN1yazPMyWCaBLu2R36jWYcmLDezyHmqdLjIDb2ugHtoJtLthP6tk0
psIotARqYGQSbY3lG7KE943k55+jsi4N9qiMJJ71Cv3++ona9u59LV1En6oK6cvGqViRqCoVXw53
FNjBnWwNdrwLrH1BEQQoEBDLhRwdIxv6YwFqTydvUXaaz0Plk0Ja5WyP+z5iHEQkFRuSmLPf1i3j
N1ztI9PYO29w/bxqRkG7kfIzvfCTJP7dtbLLRK5ozHRym00eUScOfsaK/Z//917Mk3odjj8XRc/P
jkxEmJKrWaeR3BqR9vi/koi8+8aTbP2haXzKgjNR89wOW6f7g+QzuVOWBsEgT2Anggia6AwZCRH+
qDgD7WAGKkoGyMDi9RH4TjYYIVi4kzy5xbPWFuOFzeWWscx/Ad5raUrnpJiEKytdt90hAvuRkOzc
3WQZsQ+Lx+OMl1nOuKdzeyMV0eRCGjEt9rCeedD/Y7pJKBCdHEOl06HTld0mX5ewEcc4ztyeOch4
PSB2iahgHssGQMmzl79apgKnYs4fVwK5ynDirbC4J/iQq3mMFFeRGlsmO/lfLYXEwFJ403xtBsU2
n1bsYy06h8y6kaD0iX1hvbalR4dVZnXVXhJhNisoRz5yquc56LRwJHZqx8cw3RVIgsW3rqd4Yiit
OVrE6Yfar9qsYV3gKRTlC2IgPv9Bu6+Gm+3vyxVgz30Bmn0QJJMIVuiapD2loRIsh3pbyf3qqBA5
k9gnm0ysPGoRynH9irFtTumvkNyw936HCIq5YiiG+2361NgevWoMjh+TKZrQ4aixWmyK4H1iW0HH
Eu2bzjnNmIWn3NRb8me70q6gx1+kxgkWqKGHqUfuHdJLiu3ZiI7BHSuXzY7m3QV5FUPJQDEjbLQ5
j/gJCZLqNDf8EaZntBMIlOqKseBKu9nJiuR5a43muNqcTEiZI8RpAk9yZEUnEuijKso6Q2YixdKf
Z2IEeNVulnKZyDydiJgzFkC58CqhRS4kTNAYIQwmbgQfL9D6CWRuIEvOcBUwR3KYGMma9Z7z1olO
0pRSjAfBlvA5APzfzorIYmxtjpyV6XtCmxRcuvLC5tLLEAqqjnhcd7llinkL+aNqpAzWuiWqS4gx
R2d8HAv2Wy9d8d15LZ8BZtj8QXZIUOSAuuCtutd5tlBSbeFkXxXORowvpaJKfazyrSoUUU79kjUH
EnRv81ZZi19JcZG/awKz2+gyow52QtppXMRXRHogapymHIzypYzZ3CZqVbbiGfRgNc1GAB4j4Y3k
rntWkDwwymCR2UlBB08ap7Go6s3nUCZNVWDH85tBc/63qB7GBrDK3WloR6PccQrXJ9X8/AbZTXDO
MiSj34D0avTlpoC9pcd+DaCVI8iwi96uhqgP8tgE5xn6jZow0OeqSq7B3pi0fyo4FoyDOLyTh7DJ
Pc1l6S8zGHR6J0Y0W5yOqnSRGxNX8+me6l9rUBil3n25BdpyQLSe3YYdl1XhLomwrY8AVUkFgfhr
ZE14HGaWDpQMDQCvxQxmykzAdj2se2PXmUs8EdEhbmQ/d8O7ECxRg2gyqulFf7a2/52RBPiX+Dfq
omIhQvar13nzUoYR4iayAtOc5h2RthmJfy378RrFEVkvulP4gZHgbYVYP7930Ap8Trct6UDE0IEz
MsxL/lTgIzWYXGv3zB4pFl20U2kfyBhxnuq25D6bK+330SsaqN2efVmOUbxyMoH01+GLU11VhG+C
99xrh65OYXyu/cD31tdn1Lzn9CMDIjjrCkLBOXI7bs49MhbGVwTxZDfup9/2YV1+2S3CXBkpbsIy
gULox9OPxpunU3NF3FIpDofnAfFn43fvTNTBLHi57+yUJx0SXAdwJD3jZVI41llzYS9ayGun/qRT
FdGMxY/fD9DQQUj5oAzqBgclfkmV38r3Nk+XXXKJ7RegaPdKfudYJAbKA9Bsmkyw/H/HIdcXacaN
o++vHJm+WLa4GqCi2w5d38DLA0Z5DUTBLq+Cslzq4A0m0kIN9oiGNYCrwq5DzMl5ovlpH5+nmiWf
Ly1ykfQbZmSkPsMQWkwtBOYTw70oiT10i5me9n9pnNKeli81kpEi9CISwsN0dYLaVRyDm52azdqA
gFq1QGwDH2SK6YDhG4nuQFh8d0uK+xwML4cPE1fWqjmzOCN69CbGDJhY598UTC57KGS2w9n3BQgA
B2LLO5tqESwXmOqvH3XnLzzw1iuSDqCSJMZsYcacueesu1bgBL7Wx/yuW93m7Df8fxOw81zWo30U
D7ANbA+pk1UbW4BtPtBqiergr/v0iSHEJajdvVuj7lKxVZr/6Mf7oZ3H7Zc3c2G+gI8R3XD+aBx4
Kgz8fEvzCCIC03sKe5ZxmPiiVUDhhh2AE2xWUF7AxsK6QQMntkKTdGgyAphofWGiOOLIOgkRgLE/
peZa6QIAmlGVb6rq8wm2fW6qkep0bxRiCsCSFL0IgPwFOdxr38hVxjmqwHBOdorK1JZAx3U9HzNH
k+qT4h4BlhThmtfFxEbY2oQyZSGStQCOHhqn8nIwRBQc57a0uSAs8fuM5KHMHRH4XppT9xontAru
RsdSa3gHyXIS8GBHd+XmHd4n3RCNEvMrXaeCWvE062mF24uGlwOTDT5sOvG17Fe8pKccvQ48V6yR
AkNPRIVHSoMDpEVEnUqQhKEzw/72LkfPugu/umHXSBtC2aZD/ZFOx8vovAp6qB8PVn8sK2c0tAEO
fyXKn1An2smBTCmGPbu5jmxUNDdcNrJsBsG8BT1LMJrbCd6TSiyuXPmyfk9UENqszo9Q5yPNKR6N
sxNKE6cZyG3nqeyOY6wzy68aUvRkCPMrFiT8zymsiMmCqm5iX447Cykh9AKi4UeH0UMHcPpTEuzI
UgVuVbEjNxhhnI1zLpMLUwPtORvUqAh/zB+Y8vfHpZwJbWGKU+yHrtSTwc7hUbftFKrIMEB/5iaV
/a1LkJkITi8X1nXH3HN2NJtOj2cECv5GE4BugA+eKwJftyO6xY4XQbfmY1812rcxDWWCOgbR3LFm
V+GR8if7poxdEkh9qVRBKQ4HVe6HCqmnw3KpPGEXKYf/QO0gpE0aw1QQb49sizdiisw8IfY7DqUG
3kv2so3nXC49V6XQrzB+tJOJeUWutvumAGsaQMqTcpKoyhNYn+2smerHkAGPxx6aUEfczTIg2bys
FlKmDNC1jv0lBMMjqn6y5zXLipzq4hJbZbQ8PuITBiUh6UGAI0zRJQa8KO4iXs2szDHoEYqhOj2f
9OMW4lRHhLJzB/Sm8ndQEgALiXG/RPuYnqFQ5milX2Xlf4YN5Z9xtIkDpHWq1tQ0t0H9TMOy1Elk
rngwhpLMKa7QXppDaj3E2WMdulF3b89HVlsnOaHHI0R9JCrcZIw2j1+5Gx1MMoK9ygXQAh1kCCB5
eSkAFJyXwmXXl60Ts3a0N8CPaS67pHRTLvaFhynn74No+G8jTgWIsyb+Ze1rruaqeYnPFpM2vdRy
IZUNmqtwjrAJXMuXcUs6q2TGfhva+XHLqMARCmBN9vyjEqoTeR5qsyP6DH3oRHwlvTqSLdjgqvYu
LbOrBW3AKf2AbNPTgAIZEuhnl30qZqI3NCbW0WI72RPozJChTy4JzkLm//azrBd2c/+m4hqQtPBZ
EjXaZnY1MkG8wlwucDnAjW4xVJYsEGZrVBo3Q82/UT05CGwvEC8ahhu3YhJJBRUtx7Qi/GDWcso+
C7ar+0ub/Xc6IXySYfLQaEVviNncmwXbUagDhPxe2WrJjZLAKX1oSPMxfxTSgpfXc4C46zJopHJY
pB2w0Bu4WtUhUqfYUAiQfPMA/t6jORqcS5pm7sq5MMbu/wUvMN1Xm1oUl6n3GDp0hBq52LJPAFZQ
KiVazDtUG+lqghhIqK1kVfHdsNoAKeyT2UnjoVtTqFbLEycZDIf613vubkTN0w+5Cq0LAOydFmh8
TF32/B02LhvFOe4aWFK1yXmFostEgtjvN2uTOhnyUjYbhe/xr2lg38jVh7fmql9bGt4r1DrYhhD1
xN9D5afq0WltaP5N1OU1h+RPfbGz1B1nUmFBkIG2ZJsHOzCR7laaB2StQ8zssD0Oq+hJaMdCVG2S
mv2136XS6TKDwB4Kzr2wwIw9MdkXTqEVTvaJt0e6iPLscfrOOnvOVe0cLrM+wUm12VZ92dLTPZ7T
RpVbKwXUlZmnup//cXqW6RwHl3RfMnUtGQNHHYfLQr4ENKaiiVWSvTVn7tI4JBHL1U/IjHX9SYeF
YoQZ89HMvDa4SNbue6tlV4XYNCCQqlan4fY2AKxiK44pjNSXtZmxuPfVBjtGbGhpoIHQ3d4NyoE8
7mLY/TRpUpaxHJzbO8O3prUMNM+IR3HZ6PH9uGk5ITZBdgv+PGnGFK9s8Maq5qVfdSTW2QMBXGcU
cOh0UTqy6fNrC7UyMGE92TRVJKgWeVaR6889CKBw9+GeMF8KhToKJaCqmSz0HM0n6NLuVAGdI3ia
GMKM2/6MH+jqnXabUYRg5xXrnU81x+xhKE4HumU5FU+kJVwBEckxjdV6kT0A3iC7dPbYXXrOik/r
RfIqLfW0JRut3V91vxkAnJOW01k5UkH455bSvjScBvOotLUq4tTgx4+pvh0ND7OWBrdJNdgVKhjz
WfXE0a1FzWVpc5FziuhXV5Wmkqu/SDbgj9a3XHPt3OGfu9/zE+vVksdZ42ySEUWHQ1mJq7IEa9SD
UQu9JpbGKncwAbQg0Zr9XuGhzdz8onRJyrAIhx5D1DetzQntRtzmhSlH6N5kQVdwg5dTzmtpRlRv
bY202OBHbw2cwrU9YwfuJ8rcOXSFuJKwRU/xhYrkoEKJVHSaNs1ITfP606xEicgxNZKeGgoivKq4
DP4jgYaAludGgvKJ2xyfXDtszDlPVrwQZpRS++KCCGT1KGDaw/aWUqTJrFA0h517uKNlguDXtrui
KnfIlkREZyeuD80Zjw9NdpWYLcTlWLFvjEWhTzd8wdQ18mxX73rGZq7vfbzE3p4hh76hv+P/Xf+S
a6PyzxRINuvJRzgzXqX5CbxR1wc8qRUl/tQVkkLsvZVOJ7JT7oj5mSqHeEVxlNyTaNSFt95Um8Kf
cprkYjevSNA7a7pq+JypJmw6erke5hAS6Bzy5+9Mc3R1IyBq1hp0+zSnOsIT6W6GrX2GczIWk/6B
D36EjkInZJvyIWWGhVWOtRS5ubPuWf09QxHb348kh2dZY8FBajOmA+sX4DVKbivQkAW2drALDccf
eHMgMpP4P+X3qBv/RwrMn1E3/UAS4+QezXCoZpXSeGHVO6Qe2+U0kGvtsa5HGrLGe2mbxIP0J4V7
WcAs8HtsdCGT/peioZbcJu1Inj3KN/3D9cSJ3tutMixrzD4X9HKWIdanVX1JddYwyAX/kI6zHBX9
dJ4Y5445M2995k5yXdMZ+tvm2e67fwtg+1ykI3mcsq+taKI0WZA8FldYePEwmgnAAU2qQ5YURFOI
XHCi+v/glggN3wizPLlRO9De7h+Nt/mfKdAG6guIfoJO4c0D6c84awGv1zSPWeIyfVBrUeVHUYbX
lhzUcXJtrzDfp8lm5Df1CGbhzptaWZ3remWjkgzyFFc35CD4uxdtGsDKIU5iFJFm+z12eFujULkm
XJtpRBcBtKbzid5juUe25t0JgcxI9PUzmzD9N013wrSFxQlGd81sWAODesw3M5k+Q0IICOZoN9Sz
CjZI54k2o/Uh5kxNrYJ7lSpDiPOA10WuXpC3kqZgAr0yIxKcSMRWntwIEPueNXTMgAf7+kHKcvgx
5o5ZPE4U2nIhI5ENSoECOfc3cGBjApqkLXhqv9m9OfMUV2tfge1q9dRSKEBMrJRb5nulbjcFK3qk
WcP8exLbkoVIO3mLSoylS6+LnvaqbjRM0R91L/8gFEksnaH70I4BBLns4+Trdl2RnuVPboycnsMn
Ep4jkjwMraxKBe+bgAe8QrSnV+Pvqo8FufUXB5Yjcaim66H8XZHltHl+Jw6gq0gkIkgs+57T5gQf
LMFKARq+D90C1dpmoZukrPMUcHCMvrsFLT0NFAobYdlJZfALhyzM2Iw1oscbmmnIAoNFpn/rT4/S
KpnZp0OxVlee6NAD+7C3GD4ci0K+6tYZlnff6J4vPE3u10A8ymWP6MpQgWPJgOExDSBjygYbhISH
y/AKq+bAA74hX1RvciahH01UwsyKYu/FACupjDCNHUn8bVclFtwmdVMyFS+LiTz7fQW3FvPJRno9
LTLv0/9rk2H9mfh/c6aEXIDqrhgUpRmU9J7fBSyX3+5uIZFZrtGUSaegMjms25wMXxNFGUrGuKPU
7bZtDBdlmZuvsRxaubNRIO6GiY6QV9kiRnUsLMTsUuJ0gdCtsxeevnM6FfWzn79JXysFhnDYclxv
NpFk37OQpyrzpMNRJcLZy5uVdjilMXQiPD3OckifQA00gRxWI50h7zk4hzQ/EGucRRNWH5Lox9iG
o9CD5YMMD7Cn2rEBA4eeGKezcWqD31TgxriEXktPfhJfVsHoJwTAYDdTx/+Lm/+TJhoDS7tQUbLg
eMkqY5xFGTK4eGJk//Yuaoj7bRZteut3Tb7pvN/sfoM8sq+MKz9HY3gfpsi49Vb0L4k/kpv1nRAJ
bOlJmtdDLN6XGzD3avonoivtTYxXBZDltqKXPZ6T0gy/ois/uJK92rtiklaeLaMm2Uz1lUYArwjE
C7NnAKWNIdzAXQKIeceYIIbpCTO6S/G4GzEyAmvCQCf6lLQZyWMieINYJHFr77LSvfoiPqdudNp4
A3/dfHA2VxLs3tcYqjixgylTYYxuqqktTRJ2pJoqLc8nW9HWgxMvbN40FrZSRttQYVhfX2TgaBhF
CHTSJyUktGaKyn5FXDQZbSyWyDdcS07/ny+3AqiY+tJ8pbCzrMzFT1O99yUaDD+WwYp01MlS7gOQ
5LBhJrcdwfaGN7ihxVYvNqx5jbrBSllcOBHchjzaOeF7jI1zz7NOQBS8UBgVd5DAjH3avtdNhNvF
4hhAFUx/RIaZWW4/WXoqnF8I5LJk8YRPxJODy7w29k4ao4SWBpqHOq2mjuMF5NFKa5SBOEGUZxT2
bVY/yeVtB4ybY8sD4kb1e56T302amdSI4SyBWbbLUtWix20MlV/mmNTJrgZI594+wJxpcEzg1syh
5X26gXLXQxA0q7cc0EYY0tU7pslaZDQgfRXhlbRLWy8wCGVBRIcVWKUDjRJMfz8oE9fkyEN6WNOE
jCVuin/Ihy385HqQ4GwtjQLevVgKnjas1UME9kEpQqbJG1T/BqIyt03soExNigHOIaXWg7slm4T/
IynHkr8StM5lJQm6mxAQCC+z2UCJiGa84AvBot7tq6Ypv6hMH0bBAT9hvoxFnmccnF97/kYaAaW6
XAOrkD8AmjaI/m3SXPH5ZuQPIRGE5josV5P2j0THT1XHai7i3nVvYj30RLofAEXdqHdkK9nqx5lP
4kBh6+v0T871kqNaG4SHoKNi0kDMmqmBDVpoQZ6xTHqCOwHUilZXDwKJjRwRhANYITw45ONvev6e
nba6Hyne2tPj8wDOb5CpH7tPGkdC0Ii6gRnH4XMz6ZhlV+63IrT4bsbTVYyY5lPmxKQ3zHcQuk9D
zXZqUMRCcPb+fIV4fQqQHOZv1uZAI8c0vOZXoEFpR76EXvKelhZjcaq97aKu4wp/fs0zmDfJH6rt
RijXhc5h//kSv7nuXBgc6yrjiFaPZf/bWp5nBwi4nISlrTMW2SYGEM3dMifIR92iNo6rl4qybDBs
iet4ESAnwrkMR2ZuI2xoJptW4bIfw1vJCfpkWql/Hlc9Qg4J8mAc+YQHcVkxc5bhYBpQq4DhbzH2
qEiBVJJvCGiNcygbf3an6m788l7ZoWZI2kRI/iKYZb+6zk5EyLEsfLq4eQ3BKY0OaP6Wmt12pffk
Jnm/cYnDkwmMW0Z5tfn8MXiIFStZk4T9UC2/XzV4n++qY4IF7Yi6a6w8L446GbGJVtMQWg8Xk0RG
xJJjbTTTK40i+Fri85Cco6gYI7hc2ubfsItk8M2IUuvgIhijXwMB/KSeWjMXbdySCevX1ZJadMfr
ykZgCkayN30mUp5Uigu3Sjwe0QtENg5Q+4ViUkFxBRhtcZB0nusnzoEpI/Wfyohn8NmwK0lWVQ0O
JWyddfjXgrLC3oDmnIGQX/TamIwC1l41UrSlYSKd4IYIe+x57onA/Lw/HwFfVwM/GvHOI/1nHJ7N
yAymEXo+pyCwNtnfDFnMGOUPPhkw4c1QRN+hNa3PjmtdMlXCOej6xohtmkYqgp/enB3oebKwGkhL
rS+7cwrgFic4HCfiGIJ7makFUOTMIMW+Vm+MyeJcCoHtvAmfKP2jm64s/WO7FZys7woxKIEls+0m
34Lq5H+siGKb1VIXfOTcZJY0FCnopPNAcPAiCQWbr/C4/mp3sc3XOKds+pBiqp9m+6j+B3edL0bt
4KLPeTnKXzeDgS68z81vwidIW55DvR9eU6MuOEV1gFyvKHb0XEuAgzuYjfz9imYc1xcoif+3nNP1
xTQMhuJi0p+drIIO3/xGsSeFINcL+Ny29drFBy7V1K7I+BLXbu6qxdvs7utWazrWyvRxRGJfzsnn
0kGaWLAYrtIl+1TvYGOQayTutNkmBPd8QYng21VySFdwHt7ve4n525fQjTWgRUcmrEuFu3MCwOQ1
mTq/PIcunrPJ+fxZ7yz8iMscdpT56CYppcFUtUE2xTvy6yUPNK81DBWKPQ2AyYq4kMPeTIu9c/jR
0Q1Wnjhk+0Xj6tGFdQRCApPiyx77WRLYdGLHcmWG12jxIZKPkz88lrlZvA6yWQ/v2qIfaNGJwcz9
lKoMYGhO2g3+9e4YiJoEk1lCenKZMaaKZbGR6RUybUwHmNBySCoI1p3IH4GwNGuRy1VGtp5fRTwX
J1NxA/R80xBm147H6SnYOGky05bQloBbQeyZhMvVPjD/PPVsK172qn0hYI9Yzdlt+WM2OYypL6HM
StkgHIgP71IEFTE6qwj2n7eT+A2i5a/vRosAYnwYShz+S36jWvvlPquFOu5AKFVy+1IoFudxZMe5
dI8HmA19ssjKUVM3yh0biz8jzxOIzUJl6cdO1X+ipnEL+qRu2FlinUGxXM/yt5oIgIxDQ9WFTtIQ
M2t4/WgVrcHQwfQArOIDwXDPENv2fc5P8Z4vZZPjTYtxjbGYWD1XpLDYbjviWwS6P4bmO8SV+7f4
o8SrzqqYyRj1sMXW+7HucWcFk98ZuxbedQYEH2l4czMvWnTHBBpvGvYJjSPEGB7EvSKSsmujgbfc
18hSFcF5/xRHTsSW1bBwgjGBpGtw99SfmDtTkFNNqH/lDg0Hs0Ks0UUZiXo6hU40iU2ll1FNcfrE
NXbi9FGHgyoT3mFsj3qTkovlM8v55ir3Z4FyTbOI2F8VEK88ZfJ8HNGPVI8m2KixNAATj3PZm4iu
1AXGGOlXelkwoRsSZd/hC0vtdgf0dw3NmWiZoLP77mD9+jsCXY8BdXuivNFp+8w61lSniC2S3I4n
BqlsVOkCm1Pzn+Vk4dSJpd8O1vlZ1n76ysUwL7BSCIJjyWQhkby/whgVKDXJQ4b84MAJRaPeuMoC
K2B3cEjfCw5Hbu4ytEjif95tqGHmsrya2w0PZv5dENXT596mdfRe3vxeqN7s3hSs5sC1gJYrBcF3
HsUhxUEuQmk604KesIeO2nTARq0xZJkmxCqFABWs3wODDHKp2lNqa36UKRiY0eAo3ojBu0j8LN5Z
KoeWgwQqCgDa8dxVmf23OpT+N7nv2Znfp//vFMvWZVyAV9xCOO799agwRIZTd/hCaz5rHlA2+Ol8
bIwzNCdNqrc69+RsoY5CgBGN13bE8w5DwgBfoBxiLku/AJ7tHvDUkPcEcF1FVe35CeYg69Ek5d8c
IwjMx0m3ZR7O0oSCWKQNI++59tyNcCG6PgOHKsqCB3as3s/liptlGyNTSbiQ+jhFlnHfrYsXPzUm
THKFOzyayDtxO5omFHUQ5oOage+Db9htVpZgZz3uKTKeTFB3QWNU5QcIM9nRChbjvhRNfFdOfsvY
tZV87WIPJAf5VJ6B+FRHKCe0kv6VHQFdmC1M1nW6n3eY3b7vZ9jC5p26ZEsXF2Be3hzy8lt4iIXt
l5NWVIxeFM9ELOnfZzMZlaNjftvIhR0rJkP9ggFA7wPnKIzDkEuIXqUSRA2oTtkjBb8R1UIvgblY
1/2BEWaqITRutsOhMvdj+gQqTeK2wWQZTT5nlM55S01OqcuqSGnMS65so1hBq6TPM9cSUUexUnH+
vDTxyBvvhnZWgM7I5Qpx7N3PzGs49WbGRVRoD1ixSlp1Ki9FhtDDk+8s33pl2uBGauTBno+CCDlV
KGxhVGmIISI4uHwUS6cR1jdTOV3VNKqYc2orf34PP2P0O5DXeGxx7uc1AXwoFCU8vT3naOSr8XMK
JPnFOMNpQQxEKVhnsSnEWd3Fz0E268NM7qDIIZLmgi9PXr+X55JjQ+ubZza7sfAQpBo270eNkczW
tLqm6KuLVGbOjpt55gwaJNOD7EFirNJEEXcUOdNZD8iKTT9rjCA8I01OisqHXUKoie/Omy+PpcnI
HDHtvKPe0ixjaDeRfcakiFox2d1buUwHdgr4+sN2yFF8UxdrkVAWxi5RNXjBjesbEAUfvMOdVDuc
Sjux38PzW8u7FrIS5/OZ2294AdGmPnrbhXgTVI7yL6fo0lY2j3Adws/ccXoOcRPnUT5j2/EM1+VQ
dnXc1Wyga6sGUTAebZyiCQxGqHCqRW6uFaPXwmsHfblFu44dvQ3TJAoxYdHNlmUfXkVb7xtM8jRM
34hwHGD4i97dnEysFTPP3N0mrW7qngHBXWMrqxFBs1rCfK9OJfVbVwjj72cYrhRlfvYvtRwfAkbn
dAixuJceM9/N9sVh2F11iSOznsKvvdiMm9Cj69FrBFul4m8n7BrrQ2YJ1S7uliWmb9f8wvs9Jcdd
ZY9yGcgXvlQTlVIihKbkK7+ngc4mZ1x+yKskBqCye5gFUsKkMgARtKJkpLmijIoTlxfzeUCsflzJ
WCHujoXT2c770eKSX6JC8W/pHsYjCK+JVFhYVUyPGRamofJ25j4Sx3NDROWfp/USghrL8TQ+if6N
jQW7XD+Pa2LZkydR5mNLaF5iiQ7zg5XhTM2VvFHcvIUwghSk0UeYjkHvzDMfrIjzqHDkvJItbded
7pJiuxEU1ZuovR4xQxT3FqG4FH9NycAs8DYki7Pfz5CtkRieYt8634n2N5pxYpUCz9JFWRtnxN5j
KdR1HkhYUHpEiMHOYwnhZ83gHQY4z4grmuXtt9Pn9gTM4eQGP/83ewtgz8HYcxrpYfasD4w9BpT+
X8IKKpMwe5Lb8YYeJ4V4MP0pSoYQe4sZPcvGietvWI1QceVOBmAydVcVxEAh17zM4MqIABgR6mE9
ApeFWJIuqD4ECjAgbb352KqlctVKh+50fXUbVAr//0hhX9lmALygLYxpjx82H9e3BAzH9l93yIuX
ROy9ZP3UmnEijfyJV+p1pD7cDcs70lLYgHbIViWwNsy8K4q6YFvSn2aITdMeDENCPkuiqR8gTyHz
PDfsoDeIlPkU1uYx0oAHCTVG26nmDMCc4WyhYiactUmKVhs/cvOt5zNx1nUBZeGDM+Q2dPv4su9s
q4iuQ6P5RlWyPwVXc2KfbWrhISkSkU+bMSacErx3RhTJ1xNKWLAbfOP3WEhStqp9PE5icY5pQb/0
CQfM/94zanI3I6ZYdPieClfWZVGb2NnH7dacoEDwwDuOh3x+FpMwTQ69F/haLOlhBeG9e3ZyiRFl
FlnLjRrY59nzLAiN5canyvM5fPDu6lxSVC3B+obtPV2f/6BIjQCcMrprjbyBYvpf9oHcpsAx/nXj
Vr7x7b3kJOj2Bmj1urzlR0+0p2r6VJgM6sqnBKm17BuRiYHzUxNhwgC5QMqfMEpMRWB5FDqZuxSH
XAaEHcDwS8Bxrjt3AYiMBeqq4XBCuG0CESIIozDNkhbhvWiwPciw12FTZV22wapyWcJioas8QFEU
5pWeRJBndwhjxbItLKSdWZbpcfFqVuNRZJNIi3EkQw0iX0LM7Sp4kaf5VV7nMrRXoZLhT8LVmykA
XlmKTxrZevo6UsZ68SZlM9hf/5n0qDUwAqEHyg9ckZcdg+O8rrCSd/8jXIgE6mBY71mZ2vaOX8Q8
t6t8f3T62aZmPMLEtYpbDn9RzaFmvnjrVaxos8QK0/mB+kDBwz+XPaDHT99t7jkT8Uo+ispGccqQ
nyBbRRJri41DAHI5i3gPMVWUJ2jq7mgYDzisuDFZIKM8djsA9WvOE3w8r/pY6QPiQkU5clVL9rvA
3OW71TYKbCf7WScKi8f2mLjaSRC5mULz0l65EjgutHFfPg/q+Z46ZtwKmDcovnSJlajiReiVPLL0
Ik7mGbTYjc8goIZKRrbCV0xxM0DQKZKtYltNq1WGzpopU0m2IyXFMi2qr25MzDVZNEb6UDH4j/BE
h/wlcxNK5p71fr/gX0R5NXnZBrK2dkcuJNsD7ArK5isnyyDGcBeYXu+mXQi4Qp8xD74W9s6N0K1P
L/3Brc7o6M6X7vUs4UZO9Ka6GqqwiJzRS4k5uFj9NVaqo7BeqY5r0aiVkD6ElarjFcWCXeB8Km0h
6D17BBBfH4u1yXZ+kJJhJxnRYg0QwBW9CdUdVg9bHuJ2d7PyjExJNyajn/gKiDZ0jgeUbKq6R5dM
BhsoFIhnfbese3Q34eZFRgKS+q4XzWPipY4Fdpl7KKIuWD+6dmD/B9wGZrgtlvGKfwnGDWKyKQqM
8/R1E79meSQUBjAvme57aTdg3bSo246wMDD6VukOPUmvRhaJPQfP0rDQxGHTHOtCCiei0/3R1Uh9
AYa9EsLvP3lvGoxEqTsetLVWrujLNgJSW1QBu8ik9WLg46neEYg7Mnz92S+eSNSWbwrcp2Na26Wv
Wi08k6rGVy5xR6nOybX2aZVg1wrrDjJerL+XVyiohqoQZqfck83kTpm8Ya08L7Ww18yIslS5VTJa
xbyyIjVJdVkrMXg92uEbSFuCbAxg21YBPr0LrpEPdSFpbIyGqjJZ98Dy7jcUkiCnWOAUW08QOxue
HHPLyyaHG/8h12Vcb480VO72LU2KsNcWUmQvPm+YZayhdhbmJIWfYaen80ttQQdAbiNb/4PjohE2
IXxJgtUmR9gbhphcOH4lnlg6ZdXUE+lSZeL9cwojrv5QAY6r4a0ZEr2ebbrZwv9YFyo5BSPlnYto
98oG1jZH2RIm7JyJERrCCsaskzuNdv3Vc1mq0RY/yMF2Z4REIo2c070RLZAeGwMrsVBsWC00vOo9
J1tcM7UTHnY1hS25A2eCtTIV+vXlfiiG94rpjT3/U4iPV0sHT7IkcRCjz3Ur5An4Ew9KO53w102q
d+8BzFZYbKbAx7pnMyKJ3+zlgdB8e9UwqK1w+AZink8axmeaKvPxFvpoXCACqZ79bAeKqhp8rPx5
StvQXa7KDrjMlHDHJCdwnKxt6QJcWPW5aGdFDvlLSQNv6MZYjkSYmL07JGolj+3vn0Ha3t/elVP0
UQGOCxKkJs1dXA7sfy4S9h7JklNyjVwN6DQEFBzbpT0icu/4d6C9OViSFoAplqT4FS/2EPgmmAth
2rTVvao9bj7tgx/bOaYVW8SgJt2scVLLSUgyFQsc/+4zsaA7X1N1MyV0vX/l6NAKqIV5hzHhqLS1
sm8gPG975efyjmte3HAD1QjtC8VgmNPsAiCwxe7XnpEDzSiDyP9knRcQHv7GqT2ap4JoVBo9ehJY
Jks2CY01xNqIljUFbgj4XGokH/DkNPTfFRK57TmwYXnUtH7zZmO4xOBCRgTAijvtyReFaGEvv0Xv
fgHafx5Rm+hThN74O8QmFE5yYpOMrKAc1etOSrM93DAymyWJk0h10rxmR3IlIknJaD1eAmGXXT3v
uc6XQilnouJdeKqWZJzagnrR0q/rU0E6rdiG3KTuwMh8T+qdN5Q3JZjXnJLvjAooA4+SCloHrFuW
beor+gPWC7hn8YYgx/rTnsLwtYJmiUDHz7ceJYt0M7LJDasrNbFpQwtnwuPfvsdT61IJbEb9PTZK
vE3vN3g006xkFhFInLglu5cMn4qkSbHUdG41TX61+eyeY2ewLQiSE3/B/7xa8ia1+N4ZJRb9vRR1
qBHmdWZM0Mm0xJ8A0K4g0PcNUh4GdoNtzi2ZUQScNWiC62lv1LVM6F8e52RXnGS5aNhCjB+GADS6
RMDZj+7IzWAb9bTUueZZaHuV36O2UJP2JtfdYtaSRiOmW+Um/k90Yhtt1kJlpSN+05G5Hqp3QPUV
LBxE7gS6CMUt2WL44LTqHLNoVBQzx99P086CLcjTFAts7Fbrifbdsj3yJ5oE+uMsF2+ah0ZzizyO
lNwioawA5GD1/liw3cNrWTDWWaU1NX9NvPnvmZpUaZMOuIBsjvLzGolkf+CoinwRKvBD8a+SNPcM
sSfak2uPA/Ws6C3HYDMffK10MyPLUvTBGufSCwDR0+7INabD05RvbUa3jak3S4ZV1ojLuJrgfF3X
vvlzgwxhWmDjklSzMwlFjBaoToKORYmi/ktmr6i63yNA08MdBmPyH8/ZM9J21y7hoQXdy6lG9cn6
Amo0SiPLaXs2051PTw26BPKv+SVJ25xMcbmuFF8fQAWonB6V2MJtYiL2uz9pGoiKt+9lac3bdyCO
Hbq+iBEjF5cNx/A3c6p+Xx9teBB8Jq7NzjobN3uW+f1jGNxc8Xo2x9lNqQGki5a2szDn0M/RHYGs
2N/aFptQKznjqvvfoyzpRFRdBE19l/OUnTPmCqXuamhbuhT0c6GTpAjlisei73vzxVAZ01dmcG7k
0yUXKbPwGWkmn2dG5pyVrlEXINrUYh/8JeTNbzn7xDrWGzdthAGUtVjq53KvtuWIvG3qCgY1P0Hd
qT8j4kyoin1xKTcTxDHIdTStN5D2GdkJyOFhBP8pSwO8L2A+sT7u4jz3mDWeVBdwAyiaJwAKCgDz
UAgUvEVsaK/9ELMhFDA+qG0Z0lyTLD+AXNGMdCBGaX6v3MBrRSkBSFl44dzmgo97eLvLrq0XY+oN
s+Rg38aUTIcM4zcOafxCEiDPWUZDHfpsfpYpjdk48OXGjH4gLvPHnA0FLpK+Pf3SftR6/oRsqL8R
lEwtGdirO89FaVZV+UBklKdFQmDXF5igQHyuz5Me7wgJuWM2u4xlbFomLamFu7dYoK3TXntjpCeF
uSFuWGxW4Fp6Q5gCOoFnTTxD8tBfbjjqmIHjN/7GdfWZLST2bIGE4M2enAgePJB4AAJTjcLVjOis
9UmUbNJ34ZIxaG8YCQB4dU4b1EFNjY/+t/zYAlYadyUIQbM+zIYsr3tiR4cv87lQrn8+bPUugkGu
4yG10UgK0QL9H8tkb5peAJBAGCCPGe/c2zgga1RW24kHrnou0Oe6sKg2uTuOP1AlqVpbzKj1zuF6
COQCYSgdGVFOAHFxWktL9KQyp0RcpHGvpdZG2A56TS1ksgVHNlzQzhZ7HgJVgTW/FvBp3lu90ASX
s7ZH73diA+hbimCtK9sVFrpwyf7o5MNYYo5j8sdlBx6gp+NPftc07RQ+X9N7GI9Tc9yKCCzFOJvL
Zcn/TEkG79TUUH3r7Il9dn74VuR6XfFQBhIdOYCC2No4vCACJ4H/BuelRKJCx37Q6sl+igC0Osef
CV9us8S+8zvaXfhp25sP9FgMqmEjByAt2gClyBvqAFx2EvA332AqK/1uPhtjZ5r50QteCUktmOlQ
CpSf136iRcMrQalrYKxJ2gcz2Tct0fzE+UqucXVLgtmTP9XHkJAw8wgI/gkgoReaqlwrUoR3lJ45
yAsEiYlFf4EhBuxS6XWXXGSuM5PL1FcyKBn7A8PpTX6CsBmVSVffJ2SSL2T3kIsICBiC/rP/DSE9
5IGU4cONwPb5V7zw/z28jTGCW1QnAaqK7sshhPvVOjJFj3H4k764Kab92IEHF5nGGa+i9RBnOvbE
5rEqOsl7P9FYHEbHY4BNZZ6vL5a6dlKX0rYQd1kuD8YCAF3DcUKmXcD8lIyPS/p326Rmn+luqJ/n
c0lrvb5+KOQsKRSYQ3gDY+Tw8SbtKNapmsMbxPBaq+eMlLnByvlczYFGxSuSXu4rgwcZnRW/F0rP
OuAZNZmeD8TdwE86lx9whSJFXKh6jvqDKur05ikwxJ6c2mPuSreKl1XTmudGEd/ds9Pq5vO+iTSd
5Ty2PfEDdUtiLQUgamIpOPlFLXhIZ5GaYB6t/TI4mNLDa1I2us0GUURP04VOkD32v4c169SKSVMn
qczDwOiUu12IL4ylXfvpIZqVhcaff9GEVblz9Q9NlgwydplzIYAPkuXbxmqTcgvO7ICNWYRdc6R2
h6lBlzvZYCJ+40A7Pv8BAB7ANzvnf4oMyeB5QIpmsml3hZhGo5vy4XcNZmR5hQE3mlxdTYgRv09Q
Iv75CPOploNntnWVNtFAPlAiqqg+dxShdRWTOFBmPw9w/xSc4iXBho03rUHjhuRRaR432/JTrSbu
yAsbKcD/YtqywTBASPL5MgaJ5SmdzC5e3aWxJsZrPGi1pX5iyoXukqmUmb0um4RWg5Rob1tlYC6l
BUwAbMNCjzaNJJw0sjcwmFEYkxV+petAUzb5OocfepI5iCV70ZLd5H7MBkYwuPERV2uElKXdTtlJ
r/PD7oENmevfkP102D7gg/X5emUb4H6F/XkS0tJ296yfwsA/81QF3mQhULfo6oVxxaBQ7AW7FEAS
eiJJ2F4d9LoqYfDKLKAbSm7k4+Ozc9Uv7Fl93hHhhr/qWPdy/1uai+OAvCP4QSQQg5k+oZ/Gh9N9
p6XTiQ1y9OEarm2rohmJk5kbR2GbRV34O75eSrYUYHhHNVjTFAqDXHOi/CVAagi1lQVHs62pK34L
VdI157Bm0t68ErDRrUvdMnWrleHpbnJrVNXK0aBmX1WP5Co6qdBZ+BvmSRB/33U1I7dAD15fpAi7
S+156TPqeF/oJxy8424GKycC20i9wWgaUUxdBYt7k5Rdzyl3fLKklLU0KLes0Y4GK56UZB8wCW0E
nF+XJw+HA58SO/cnhhSrC6KWiK9QLDH4etVUFTo5yKQ0RpSC6lxuftL7fNDecfeWDvIJi6sXnWC3
Ti6KYxNGk2HP00vDgnDWfg8LmRrFTH91AbbAKYGP3i+YEWDJJaByYK42TJJAqWIiMl+51N5diDV1
wdNLg9hJGeFO6LGJwpeBnov4LkH8/eUG24z2TRbixlPlnNtgbQAoYKyLvUKIXwjabb7ZOhk0ztvQ
4KYBn/it+d3yrglytXluX2ABtEU+yKoPwxaurfRjpDGcv1mEvlVI5ygDr63E5qv74tqHV4L1Qhq3
UhFWGyk61FTpiw0mV3DkCTE9xhImtWNo5yhgtDigFnoeAsJanvJirqQLs40gzjsOETuNtSM4sibk
SO4EdHrbJ54q6V6xfmTx2xOxKsAZBXjqeCZk4NA1rOqUf2HeEeqwwqfSB8qGtogT7sv4aoJHQdzt
5xL6iKJnKH5t3Zq4zzUPAay3QGp3Rvqr4VhVTY5qK7bxeq0eEih0YWzkHGngfG9j/0T76mnB8V9d
dH6CRpozmfTQLYvC8sajNCfL6gRLTMObPe13OVsj0HMk4t1bnqMYXauKcxCsIos65f9Utsh6hueQ
w5r7+RvdoqXwZa2zBPPkf4GmJUbLlEMAaeO6MipwB+/voywzCMBHAmVdKNIhWwD/+9ASX1iC7AYS
O90sOmdatzRqiqCb22ntWnhZRJTDTQs/4jpiYo8GvLdt9xRd7P2gqF4FB/lfMQW5kMpCUuUyr2VF
QVJ50ndEkETbpGbazfso4HUJgTWIPLzkW+gEWE/CX0dDymAlBOM7x2uYHMfxhJiidPVF5PIt6FWD
tqhxtUKx25GFe8IEspUjP8LmwFNpNV5bWrDt/I40INv7C6KvmDqhbnQNzYxCTBm49CzJnkLaW8yw
LhcexAXeXNtblWZh6l/iFtunfX6+SVvHWTU7z/EJ1EZ1CAJ5nDpFQ6M4LAOdft3VJZOj8Fu84GOH
lVGM2twd4LkFd6DQJxPqXS5jme+PtMV9fk8gH+Pf4YkST8+DYw70kneHeaV8UlXv1GLYW6Y+sntf
JRexKK114peS0htRdvSPcU+ea0gAWGUkw2dE5ntRIKAGLPbHuq4qMLzaiPndo6CLjIIKEa1DoZec
nVT9g8JEKwJcsIho6eqW3KEbypTtTpi32QSA3+Fq/7osFlC5vWt9QhKuhaKyCVD/WTWVzGHDVmNv
hrHQgNO6fZMzZKIVwpgPQ7JRdKhMseZQtxSqYQiY5RIR2BlWvdAgx0cvq3jzqOzxObvv1DE6/3bq
wGpfOvU9u2T9YjJURf8FdlewKkgzspMeGpESsd2UWsePFcZLcdz/YtaJB3Qln7S2J2O4RXHx8rU9
gxC8L00H/qz58KuQRp/fKNZpT5CtTHTMQQFcb6E8j6955fA+hueTOBhNJJ/cOre4sQWPXJiiLShc
fcA7PdCAbbrYHEPl3N57HJhGI6ivHqirzZm0dxE9rYH3dKocea+yESkn8UV0F/AsLBLkncy8+xW3
mgHhBt0Pe9fCJHZ9m6Ch/ctsa8eOTEoAhY9TcbXTPjAFbwbW9oWxR1lbCFZkYtZ6zm407dNm4TUW
Yb7dGNk29v6qtbqVorww55BThGSl0CYJ8I/+3JTBsELS4o1YOIZ07WTuZZJIAaPzVCw4lXBQ5Lgx
bxdf9oD+egCnA7/fpUY0qrrm09gubS+g654mNHsFWHtic7ybmWhwB1LnRtm+Ej53iqpwb7j54HqL
1CfPnEwRtXdSOQy8PMyt6+cg1WlI7UUPXZmfQLaPNpYatXFoNgg7Ymz/7uJFmiMAgn7oLxPaEISJ
y4lpf8i0y+UC0DMIxT69A8R4pfuHqI1PtMq3JJhOE6iufBaueK08UAexBfE6sx2QRZ9+/B2fkNDB
T0iGgTV5IZZ/zgI2t0RoElEIW6oFNmK6yTVAw6gtOVWx2L+XCOIRFJROE0lTrfl85JhATzmhOcV+
4ADimTZUHCc/Lh8ARY69EGqi1uTq7UdV6tgSj0fbAUnZGz+XPozFc3r21bA39vgBkMdnrdA/5T/j
fBaEeW1q9is4d5v6H1JSAC2cxs4fX1kr7cb4wwiCDvCCXi859HbWZlyM2NKKEJ0K7Qfvd9B6Zzvn
vED9BzusIQz2T5CmA/kXoNuz3rlbiyaT8tLmjBr3NBrx78ve2pvkiNC6iDG46BAIyEgTK/txt1vy
MzdmaCSK/qVJVq/wFdaZ8cabohcs9ALT4JZKOPLb2cIzDwOaekaKCYZx/5/Z5uoUJM99sQxw1acO
qRPiLrIU0k2KcvIEzZFfpenLTseLKk8bI8hym7ybFXPZLCSbh/2UKYseCU8htOWjKVZDdzEQYDmc
cEf0EsheFrU9BXqUbtR/ENsDKv1ExRFZGXS/bxPZfzLXH+vqHzvbp4e/GvOb7c4Py6OJO0Ver/Ov
LMhZA4WAA1Lcx+CGRQo4/jcl0MruE4nSjEcbC9ILwTV6jl5ukf6VacRvxyhXdy6dn+KOMhh97NXa
njURtEo0LoEnbRro+URaq9q0kiLD4lpQDzP68YqSnwqbAg16w33ImvjeCVkQy9ASkALJTIcGoXb5
NYXY09DInyECxx2fxb/jJRQdmN4s5F5C3q0StCj1UGL+800lRyhBFuFo1Anf1Xv60thR4uftUaT+
bPro9sMwJOTbGYmwOo1RsdxqKUtWYDwNXyQUofcoEyw8wg9UMxfqjlykU6o2WLSyzhJ3NyXuCYFf
qE9qiP6ScbfXoJlyZCrPm0qZ6oGpB+5NETqtnceIpgsjoq01+/dXJCn/aZn5PaHQHCV4iHcXeXWJ
qqkLXisz3S7Z2MXBOhrfysvhPazE6Ig8pMNRDkWuS/k/lga8mpy2gz3N2i4gkXC6zd3Q4D5eiyg1
omJKTdDS6b1mXZCvoJnxVkuJdfgEOYeVr2K+i3OmhtScAxe3vqVX2J7aBTbqkBuds9fFYN3mXku1
l6IOFJd5gWKl3ISqpiMzEYxUih07fropACs30s4yKf9LH0fzX63FYTjQQQ8DTRJAWZQQaldvfBcC
ioELdK44uvL1JViOtsYm9P2+WYHWV/D2LMBZYRgIkPpWf7JJ0BVDYmusQ4DSOknDpwSMjk0Gw+H6
SmSe9ZKUvlzBrV6kIqZq4t+mylPLC5K8ZOwmXq0N15GKldHJLFzs/E8nk4FC+trBn268FdcwqlDF
sXSa4BGCw6ZESPztpQqaDvJmVxt9AO3DEOI7b5podeTOBcQiXx4vJCQybImtbx4Xx7yJgHN7nC9a
QOtQ0ZjbmGXDZ6uOXaeKUI1+WV9v8ZJygnZlQ8TXLfe5D86BzU79Q9fRUDHv1IgizH1N/4c1vf+z
vVfEM4svvjTC3yBj3dsSW0/lKEy0HrlXReDK/FfVhHTRIZbbTpNV6Xxnn+e1UR/OEWm/3U3dCwAg
tpGXp4qOzDBcDPryl9NAAmquVUbi3UpuXG52W/nTQHdyFNY07vtl+Wo4q4iPyiapA2k9KVXLs/2n
bOM39hZH4j6zdsnW2s4Bea/qCpGRo4K4z1TvmpyfgWDiTfFJfEE/eT0YAw4RYVZC0CxVgfRw2Ngd
mvYFLxZntSF4QWkVWdGJmS2srDE00GnI7ziD9au6fT8TY0JrrFU43zHrKmOTF6uEu+CY94cugdDm
8EykUXeGI57BN0RR3luS13C82u4ojBOY8saE/lFEXHutxgrAIwQKJ678llYMZ+slOvOwzUQ3MJwB
Ctj2bPqjuuwyY7Q3gHzTO348LX102awDHKIBv5sp0kpP4wnEgG96QLrQNDLt9bHUHf3RZlh3zGIC
VL8OctfQ+PTqQktQ8u76Eng+eR3xNS4WPhL9I1AJN7Nu20TdZjl5Avqp3m31TWmKi01jueY8EviR
pp1Y3/CSwGKPnYXvM0pNtLFTPtElFCzzEtlT4z5Cx1XY9oFVMVsmeZ1W1UKAWDPhuh6UbXKept1M
9YnEjcyjB3lN21LSFMCy2H0X9zOH/l2xMXKc7OvowLVppIIPq0sbbOvSjRqbsqLHZkQSyV4WVuv7
7tDskPa27Z76wl03OktRkpZSVKvpmPQYnCoFVdfddAb/+aZkBkE6LOqVM2ASLd2ejCXlWRcaiLAx
xj1W1DAX2VvRqClAIrEZsMHHEMyYJf80dWju7sDG/6y4RXRLhFm2+AWUDy1DllfoCd0WcnYpwsme
LBZOifHd/VzT2x8CBJflDXB6CRlamG9Z+eke7TrlAmfMFKDKDAIpfwLDqX8rfmV+MaZgcDziP0/f
TR7hfGyRvgCekICuctpIE9F1FIcwKrJXvxSt2/YiPO0XAvTcSddL6p47txYhud1tmeiFygrNEIqC
SH12WEm1ChDCByYmgJcNBxSYmOLVUGr6qcdwWEOVkydsFN2PbjmZYkiTeBTI+ia6Kr9Cx5xfNR8O
2RotQAN4SrWQFBIMHQQIxFeunJskOz2RUv/3fx2jMCAkm2LOQ9y+tqUJuoCcGwS8jWgaEVfKZZXF
9qZVIZMYNHkJ9XJuxV2HQJJEDp/B8lThbfZVDFaJ3aARAICsz/19VvfMTB2gD7yNs//Jo/sCscLa
WYzYKGnaAABwakMzQ4MKRciEvWA1weD48G3YHTUwxyYUniEv5uEd8Pyh53ZOQDJF+a4hVQlacQWJ
F6rET7jyJmJ/BGULccwkb3oDoKPL9+3WNUCzcJ8aPfzvvCriKm4XgMmTrEzVzFex/R68qDdXtz3/
3bRAPPRJzE76h6TX+2kIWRxHGJeC6esX07DvWsffB2Ku2qHsaMCmwDh8wTodrkRp6x8cErtQU7OU
0+BeAIc23ARoNAwdiNpPna2XnPpcjM6ivrtF18iXWYGTRdjp6Xs6xsvV1UdgPp4RV4YF7FApavEH
sI1VZbOfjCAFMJaCmZHmnC/5BO0hTW9L88m7bdeTZZS4qaMm2ZTqpLg+4HpYYdXtiCLDY2fqTRqb
rF0a2ngGbdlrDvaGKVs0m0ICk4tDSSbj92oxBIxVWsxARQMaOR3vG+bi/eDQpNWPHVElusrgNZFR
3YuVDwoyvvc+HUE3C/7OapXnM60gytCwVKUpIapLW7vxRGDWpODGgad/pjz/0BJTeew4mzyN5XYe
7DL4+qbIwBgJExYAHI6GYQ67eerldFcd0W/UXjuN3/gI6vSGgkf/dEyJlgOj2qQ4ObjN6TVeCu4h
xeSkoB59AGT9AloEiC2QN8rgpFG0I47jQt8xRq0P2EMxrLXyNw7hAQ3AhK8rFCMpwqY2c8Pvuglh
D6xCwEWv1W/zn+2lmzKcvLPEGxvUudQBLurXP4524TqCuuTeX86Rpng73uK0NIyYqr0/QdW68r7G
8vK/EdYvFe6VT5WscyuoeyQJSkrQhBL6y/I0424wNX3V8YCVxbnFBBTnLMCEeVLK6cf5kJUImuj6
vfuQndzJe66508NF2lD3W4VBtqVqDbpXTEts60HWRtRqumYATYdHWwZCliubWDPzmSE27RnHkQTa
eTE93QZNUa2yUEJn9LAx1xbB3n3wShhNAiJbur0gewR3Q51fRjpBqMBKQB7RheC7v4DSICCBT1Qe
m9ZIGWyfeQahfYfjP96QtnbLhvkrm7H9iWGsS34poO3DtGTTQXEs648fLpN1Mg23msZpkFc3i5tU
2bC3nkLQ3oGl6DU49G18VsQvTNtVH/oaMsAD+v8ZCHKZD/29AWKJNV+U3hb+JbCCQZz8QNcCrnIB
I7U8daZXw365+Pl8UfX9v6GyWVwXFlMu/O16YbIGz5PcxkVuyd0dpE4mLu9GA/V35Q2LNqIBT+3E
UjYqcx5qUQoQ2caRaBcQP3/P0+2ouuGzbZ9+Sft0igLnKjQaivCazsQDypYhbmez3y6G8MeeMFso
pqmDQewbVM+g0ERBby7ismA6dmlY3gctJgDYrQoqq7WaYSp71Xv++InqRmpuDtd2ujhILeFr2Ewe
mPzgLb+4XoOqSRXY47JsAdlYugpbyuoR5A+yW9xIG1wLi2tQmw9SArIZMsL/EaY+z0WyQ5rUIvCm
0Anm9u0Bgls9Padsx3CzPa25HhhDBgCV1ujfHHS39cpqfTb0OSbKNg44/B+Ut/UQS+hXYpFtXwPZ
T7nKwAQEWIy/VucoMyEiYVspz5iJIZ3ytipfnjoH7dgaPR9LJ4DOM7dTzdM9S7SBmedJEkkrxyUu
w43qJCvX4eUnlAoCzHI0Dj97rbMUs8U9tku14zPccJsVjvYEaqYPxmhfOR+Q+Smj99NvBsx33+mL
qJjiB8z7GxdfXrYn0XtV1H7DOODTcTrfA9z2CXxyAYq7aaXq12R4qst0/M+VedEgR2C5oXfS/Nbl
H1XVo8DwKAojNUaEqrD5WNyaacBTkRDhurhEkw06SBpnckpq3nC9bFO3ekE0O4rz42Lg0p7R/6ih
04RQ3m0ZnA3xMJJOrtDKfSxyKgKaK5LrS/lyY/lvhdEP3l4lmJfFN0FLnHaVF2/uIFw1V1Cwsswv
ZWvHVOFqVfxvk5wjMH6sU7g0pf/fxBS8p2JI8CW9i/tUacUXDewjHrMp+c0njCC5jrBai4cu/ZYa
QJMU0ZlxGPhhwBTqJZVfi87TydbXOJ/JUtcIuDv8hoAzMYKwhz8hnTcUO3F8ApUGTnKaDswpHmpr
fkbMUwfuQ846i8E65D4w4JFJrJXhzDtnAneeEdZ8nR8F6srrYT+rDzqOC0f48GWhkMhqLWUjPzzV
sDrcpsgkLBH2gSjWCJa8dHbShGgX5qj7cTxjwYeWeP3bjtsw7mfgje98ZtLncl3NkUur+MHYMlTC
gdYbP5wzQCKLlDoMy+xMM6x0OjCPYL7DRAffPL14nr3Nnd5riK00Yjzn4zcA73vKVfj2juvKWsGZ
A6sQTdWYSxf3aLTWumAPtYO4ctm5xbbktjEakBC90SdKHbBLN+0ewhm2W5eTucn8Cp8OP7gzb0Br
IdFI0NT/ZGprjNn9OfRtxqJW0LZ9BGX/AiYCUZH3tgY1AG9ZJWcPunv/m8kxOTKMahLRJS5pQIRE
iuHX7p+uqkU+Ej/HB0bhJFXHBTxi8u4XNFlafZ4OB09BmulhT1xKEuX1HtlN+aeSEzX6n1oZpX02
oUmfp3HaLsi0TL+9S7ZC1QWJ6UGhBNrcYhYfbPnWVUFXc8xONWTB1X5GHbpUqtGg3KjBJY+jEKkI
c72aIcXNSXMka5xJFmamfTLO6q9gIuXJnh9tfVHfyOsT5deqrQBbvrIb5GM88c0WnnSJvy+kETjQ
wfvU5Hf4bEmHwPTKkNVXr6jOnWrHJDbywC40w83y7YNELaS7WOyt2bZCiGEVdjh3Gzb7PQ2Py9eu
xnlLGh80i88aBM5fiHsiKUPeFjhG0MHvryX5lBnMtNga9TpAvtVr6d36PVuyzEqIfHhNH92dF6JD
V4huStn1rjhCM77S361kDx6aJjuwFomh/B6euQ3Wg5ZNFFPGWOgbU6c1jnom3rAcixnIPHvwfLGR
D3O3UsscI9aapcN0hKdckbhG91FEIMGkcCvVMMJcbPBmRlSFG5Iu0R0sPDyVK/x7/9m9e0ITEFvo
0/dn3Oo5ND9cfR7Gc6KgrI7k8ApCOeRFqeqZt6F6NfJ/u0ROCgzDIkuCTph19rcsblkM6DR4TVxt
kuJYOEkMEOACEmyonQPF7yNIKQo35tPK3LGsEV/pBHBzdLvmR+FxMjPPSIGiJC69NXNXL16OXS7K
oYRZxoCO3XZBzewg9aS3WxfsJ38m35lMaWlT/tybor/UmEt6Qw6EsZA4FKLAQx91kWoUfP0ZuyGI
/f0+xNVmlYf6nkom8QsBQI3HHdqY9Mh0BPehFY9ZWS+n7wg10FStTp8Ka/dUihPwfewlyn1UOpVB
jfQr00mh9dWSB3Vd9aFAkRgaojdtFB+dhrSs9EsuqI/JtaxDYKT7ghwcKfjGrPpEbcYf8rXx43Th
ej1EkZQ+qm7IYD6528BuU6SQSSSDFuwiYbvbXVqlmPBlxaaqMawxpENjMPUuUTGSKK+Xln5a7kvB
IKd+L++DGacefXWyH/YaS0M/MwPy4nLisa+spx4XLtFN4f/5+p0xXROG5V0L8fqS7gw81YCUsZmW
FQVcytWaQslZ7y0xGGqukcGFf1GF6gY8PAAd3l0PWxx5jLO4TU1tENsEGeSh4mEqxlE3gIcWD1HF
3ZBUv73/B+wXz7nfOd8woWSwVfn8WpcromL5XUl7PHSYCc07syVyn3nWXMHL6uUfb68NAoMJ8Ald
Pz3AwLKmoQyalmzKbfF10GoBzeR3qRaeqJ1DyWtCOe5Tt7pqrf6r3lREBNjGZyIGGGXUVMH1GrRr
3xwWwe+1S/YP2092Kr+Hnykke8u/k96XjKnjikexf7YMW3lyqIl7WJQrgWOvo8x9KYbILGmLtRjO
4uJ097SCkm8PuPrhm7vC2Wt5ZkzRTRs3T2ObsHQ9unV+u0fFzHxyHD13Pbx1CyeXROPRB8LyHwHh
tivLPK7btHhrY4nFfQIQ8HM4Q9DR/NlAZg+MyVkvfdG0+VLOkO15IlGsj0nuOOFxqi0nHzauyjTy
KaNGpThbTmdcMyAo4ZBHgdwaoa7pTZCKYbId3RxxMX8fl6RY5oF+vpAfkoV6AThNPucKDpZc1zVU
UrJ4WPiRevHooc8HtN5bjdV5wUmuiKSrn8d9BV5Kvbz0q/or284BLgZZ4qYk7GU2/oaMqPo5fv5I
cCXofeLN3uQdWUhzUv6SroxURvvaSGQy+jqXRofrNq3IUADYf1x9jHJyaF3ssCQDYFLJl+eoJ1Ep
CioQQY9p0K/6w37L9M56D3vuR8XPZbw3XhkldQTd3rVSe5vcIx91KKVI3fZ1WpNocIhpMH6y0Rex
GGHlKw+wQFz/X2KX4iuQb3p1pCBwLLNB2I/iuk4nOloAWDqRThp63yIafEFbJq3S4+G5AEZhTlqT
epNg5bBOdA+sx1yMrGTzLTrbUgfqTIQT5qX7P8RFuwRGDDbqPZGslR12kHFwiC6IoYjniH9Jqjy4
/ntCQRyVnDMnLgK5HIitc+j8e31ypTVHPNu242LZXFO1W8g+ydiFUXisJCRvauzneb6cqHST+RGO
mfNBOYgs/Oup0XhQVnLUFOqHMpQ8fdxF307h5Ft08vY0KMAasM8gTkw+hWqAg4NeHVJCx+zexca8
KuHrWWwtVkSstHCDZoSdFY7uWQtOZjhl1EKQQcAx7nm3NzQCr2HY43VWuVhZpAl9+hSB+z4qnuwo
DbZbw2m2PW1uEZG+QQmNfoUQ+zrUQVUSy+zE1FjwNl81gLfqvPg3M9/5yCV93kMpqganu5SFvDwO
RdnqHr6Zz/vYx3hZOhxGsyaFQj4WrObIdht0CcPFYfJ8zcKJCpQ/0U+FgzdTEHZ7IHh5tK//dgJg
sclZFjmp9OFS4dIUascLSXgonvz6jG2R+xc16QZ3jGeG2ii5TkDk0ZKMQec2fF+ycYK3dyzABlaF
kae1eoqXdVhw9uIT3LH1WC1QyR2tMBTMRM3P5dojivDh8FHjfpYXVNSdes4YUZUovj7R1/zQL20r
EVkvj46Euvw4RLkKzEcbHtgM9TZ7Lk0nMqt0Z71DgGWmOSn14MQsXTlm0Hf0QpIziJrY4ci8Fg8V
/M9PMb53eI9hKQGRSFUgITnFlFAne8XsJvmzB03zmfvM2ytUBd+TZV9OwSOpJG6yIEJvUzvV/4mt
VwxAQOBUgNeFdIaCoVoY4LOHXP8tc3WLBqpki56sSWvGzqWw8GlYoTdmx9bhT5VQnDDxtbTRWnhZ
PxDoDNm+GiN+HCXnRRTpqE5WcVY+pfbLQu8WCiUwUfufG06a7EnWIN9Vh75D1+mBfyQ5bTE6EHwH
U6VM0nINKlzAScKfxgZYnTrK3Qdk8qYIKry/574FBnM2Zd4RgD4LceljiRYZgJQEp7Zx/jA+f+KJ
NgISeh25FPUHq8hysUbJ27jZQ4MTY/edl7LiFtHBCwv0UlJSceGhRat21h02Uki/RoAuKM+RuzS7
beCrm5wSBL1pajIzHS8Dpj64st24oflBOZoDf2Ic1PXih/pEZJCNbIryG+RI6R01DCkaJkurDAZd
OeyWqOvNe0pC6B1zsduRIKV3/nNcHenrRAlyhDr8Mk/Ved5XMwvQD1QkD5ybaIbBSopckvOXECW5
Ygr55V1Xh+VWjfWc1lrMP2eWY5if6SEBCnNumdbh5qLUBfDD1nVgGYlG6vLbLEOJ/U6dRQb8eJ9n
bOPRPymFxqASTAyXVdqcwRJ8A0gOkgX8pAa94H+sf0wTsQJbKz4WpivD1EGvLmN7ngwrsqJdqv0Z
tOwpAWVTxCY5gMKwk4DtwYeSanVkTOiGOE99htrlxXSE+nK2sDv00q6MdYUKRUuz9jnXSPFyRvUa
Q5F3W5xnNB2+cYQn4pzlY5qEfB74wruVWHVL9kgK+fdky6ygOw/hm9R9x2td4jSdafzrXfgDnyVc
CtDmFJ6joUuNS3jgC6JbnRtMSOnfheo5d/xL+ITS3Y2f44eEhCfx2xILgHZl7q8wKhgoH4ixyy/K
t/qJuIz+uQI2ePhoPkDspfOx0xQcrS/dAxiCyByFEANU+iOxFHNXmg6kMTZvU4UZJpW9/C9t3dWD
m2p4hcApGsJ85dtGPciIhzFDgkCCvGau+NXKKwyPyhAfkfhSLuIOWsMJpaweqsgxbVE3a8ONIAo0
BAsGgjLobfVRjXka3sx6j8RMRXg6Bpj70yjN3w2SDN/kdvrZ3OcmDXPQ5MS9xyws7EJEInB2y5qU
kVhLTtJjt2kGh+bpDWGqNSfLXzrNKfo/CYjKzuxF+EXmHxamB+32H7I9zbun+ybhPJezLrbkhPeb
qml+TSznL89oHMYqkGHOMrXV7l2vwxKUmIDmnmLAsR1jhTkcyaYxv4JXBZhKnZDrbZhvjCvwyRNZ
p6KUdgWfFiH0e/542bOnU/4Yh9OV4jqebqogHXeX7Pkm9azMiy+kH3KYvaKRuOkL6x3BnqJl2dmm
85ThYkqdhP1nXUo14NOqE++y89zovkFxOqNtPVizC1/EiBys25exPHfFyEFcUZ3YumhfgxbCtoHD
/n/fG+OQwaAwwm8wldo8QPIvbac6tG1i2lRwcLfmTYa9448SsRGiQ9CTEVBAQPTYP3IkUkOjgS4B
vuYj7JYotWv5IwPmzAfLHsYETchsn+T50oWDTl880mCvxp4QfY71ECnpEyBf5PcXE1SHfSTKWxsV
AXL0xf+mMfha/+arcqAVk7nPapVPS4zs25EIXOkFA/nOEp9Eq6wuzeD6llR5plFPTqFtCtmceu81
bFzfiURPyeYsoCtMz/8nl7CnQQ5ZMH01fQ+Nkgnr3EsEI3riXkfzEtgEgNbL8wU4UurmzNbhEYrs
OSWoeUmWeAcWbHPtYEufEyAppIwtS7Qeu9VaPK6kgTEFsrVHzRqICqMURGHy+opRQDc7/zPyF8K+
5QEr4oSp8tbGKAtY772alHq8xqjdZF6tvIvuFUzicAUf/2sk4rn3v74C+QZ580cKLQZWM060DFd0
Adu/IKGFT98XWKNsI8eo+Hl6j6nN/2kXFebWcFR0/9lhEMgCVghyG54hQQOsFNZ1J5YCXNMJxICB
kSVdUExmrHQwdogQ1WwPD3gaF8BZx1dnzdowo7N3GKzgrp3c+R5scC6Y8MiERIyZSLIhbDr1Jx4S
di4EVjORhxf4i3OsnoQbSNhZ/c1J99Z2tuV693O0bA19XIj1RPnzFeyioqRyOze1EGvM82MKtnbC
iVBZyXE54YjOADmmwmwVC9ErcRiY/23rBjPuS3ECNzyO3j9zg3hZ5iI/VG3xpBDv5A7EBgc67S7b
+iQ45ftwlrga1HkjT82/ovHha6oFjXFnOuuRoI3J1RlChTRR1bU6UcTZavaQigB+P5/1gjFQKDBm
G7EAHuEQB5VscZlCeNgQHgXFJO5PkhciP/kh8scP4mFKK05GF1bVMgoZDUNku49idRc/VT6nrOQe
rAV7HZrcibGg2ELRbnzB56aOCZ2USeAen9ABQtLvkcuGwtrxaasM2EtsJdr+vZWWxEyavbjGRM53
3pW0HcnRBeA02cMJytlMooArsE6EdCNZhmNpeTCU+uguvUvw+awuIzCbTaRudWjkbU6iQBh79wjG
K9BZz1YIcQa7znmxk4tJqqYzHUx+8VkKHtVp4uxWvzS0XVIs0OVbaV3FWMg/Y6Khl0juBhgggLnW
wb8iG2U/R/e//SQhniyTJIoS76pci56p4W4zFMCgxo6eLm8r3y/O/wm5oWofZo9DVixPtsdfWvmt
rLIgl+HYQLbIrAnB4juKtnT702X7n56hHMF6CydRa0wbFNlpHKZyBZNf8hQeK/Vc/ahWzaKm+rqB
byxGc24QOmG07NISddN3g7rU/D6M0LFySBmdiRCDHwAJm0wSS3QXJTyV+CdgBMTvu4kZnGh0+Xta
hcBth3ttWsC/0eoBBE/iSClAxuCpZUPRTGDhWVYrLmubF24UAsa7J7pYxafOHDqsu4fujR/gjYyn
VIPzDNRXM95WJeTgsofjyCiEp0hIe1W0xUmr9Ytf4BVgVDAJ8L5DT/q+xZLKPdX883gNaTW1WkTN
glLnXGgz2wuE/+0Z+eyae2daD5i0s7Ip7xWRfxn/e8tY5GX9NxUCE4MVo+x5LIz4R/3/knPz4/oB
jsSaQJd6p5Gokd1Afgm7ZCyug71ixM1jbyQWQHPkr9ynSsz5NvN1JkLHeA4PqwtGNsunL71mbtwH
V0B9lTZE7WE04FFxwnmjBrX84kkDdf40R5iUAR22txeMaOM8wMzwzjov5GXg6POfEzXRfnt9AwT9
F0FxtFliaczTnP6NDJzVbxT1D+vhZ5WhT9IrpdMge0kA/HFbEArD/pCedCLF4zmztsR16B7/okXL
fk8wKudVt+RheUjh/m78Xkni2n792DaeWYPLH5DBMciWP78dUXidLT1tMNmBHzPyj+v3roeVuxhU
jPeQoHWXwCn/lGBU7+BWz39oRTvz3en6U7y+J6le+4dM8kkim4OcxeP2RbNbQtCSQBJuagBeMtsZ
KpTRlGa0VRRNaziqgjM45QqR+p23Vfs11Xi33K1eb1IhEhPWx+eL5N4MYgFrGkYGFjdD8R9sxrq8
ew2lIDUMxrfjCDVQJdK9sA4Ow6OqGZJEwsHyAnFkA7h39/EuyA5RvbNxiI7JkdV5uR6ziHL3U9cP
2nMwEP8P7PqnpSVaudrEHxbz2OBo3Bd3YOaEA+3h8HgAJdGkwqbdGos+DgsNgCEDjb739PNMKKtj
lem10noQ9JOBCUci00Gxf0vNtvOGrb8DHsAhAMyxZq0K2T3XbyYoZQmkbkZz/Vfrd/k+45rMvVnN
vm+Pz6eXMTl8IKiHHi6JF4misudccF8J1joWWuRE75Pu+CG5f8nIfgYCXEbNP5oqcp7QodVmunRv
9r/1MZHWHqQ3dufImvMJDHy00hqAywLMtHllinL03g+LpU4x8mwts9d5ftxe/gGDXiGZkH0jyPOO
G7ybpWsWOShLzOOFxGMTGIAWRSbj6KLrC9COx2yKdlUKrwDQmH7yHccocV4aZKDevWS+3rx3JeyT
mGq+o6dfhQfE6gz+xbKak/z/4B74Ekl/XruJqej4HsFpZwq1keCBpH5b4+ORzNPHG5hvfgp9N7+w
iV9ydrCOdDl5hQw78dtKNOjyTL4tkc/tiCndTF1m1jVuvB73O7JSQDaU2ntlPn+9vhmXZugZ95hC
a2Dbr4XkJLHV9BvwgI3JXEsZhCIYsQp72oKnQP368n/EV3x4z2C1FFAsBD+9CGC8BOf8W22Fg4AU
FvGEXG8yZZgaXLBwiS5lh49zm4+eItmUTYlrsa4yVCoIyj9FilqNI1b8SPehE9/2byNweSALQhM1
TtBs9oWiv2MokRrjttESr4Y7WKgEAg8u9QsIj71BpI22hDLUM5bRRsVZAxjOJZZ+N71cHrCIzklO
G4muuIZacTwTsWwI00h4ubiyhAx0zN+ev3U2AgmtSxUV2yJnwhCdwfXP070cYTHwxFOWvDo3Gxh0
G4yE3bX1QD051jyTVdQdA0EGfQpE1wJLNYsd/g4P2PJfPtjqAYRi7jpAFBhPDhxs42baRkDDYy8w
2ikh192VD2f66ppx0Bbqqu1mGFFswkz65dsdblNcWliwHJLJ1e37ebZR5l3ARs41Ib3cIC9aVz/G
o8CitlW4XziGoAKiW1vPBr/tAt3ovlNiS3JT/qLo1a67n9tkYVCKR7a/zc5NAeDqI09DxFDVfj46
DZqmkBrNPiXiB88siywVoee4Kw2Vw77dAt35CeYYwJttVPhC3Smr3h89ou8M9cDxg/maYBj11qeB
QZEyDaUMrcnWhwTo2xuDjMBj2wrPfKYkI73Pr0g9Ao90Wts0tFXK0KJAXl6m0X7Y7juwv0fFXhd5
wITAH9iyy/405i4E/0F0ZFz2aOyNsYs3pvPcclZjau2F0UUNLzgnW8qw1G5WFIldLAEd0tIEDmkd
AoHrO/DkUFYC/1kphmFubzKB+bQywQw6cGAXMoGAaS6wM+rs/U0u2iwcpvhnTToxZ3CCeySH4nBN
jgbA8t0y7EY10zfHHNAXAGZ3xp+Lrvhg9uUriPDrKygxqfCXUbxQVU/A6Ffzmu76J0wfZpn6ZtxO
fwurgr+0CfneDRVDBfeLI63Wg3HAE4gEYTRbXm/i8i31e0ERauF57TFpkRGz/o9+c7oANgXNVytj
g5RLLuJFj2gLrx5/W6LhOAQwAIYQrx3ZXSLsMgZ43b0hsITOOjhIiSZFUGi+mBX/APVAFlmCPuGG
5ansB90/o7QydC4P651/BdGDWE3CSHE+tcxcB5Wb22NyuY3s6OTkhX4AJaeRG1grcqVH5d3TkFAu
i4cd+YNyvrWnAYWKNJs+kNUGreByNfasCADAIqsf1BXJyfHr6mAmiZVkdYpCv2fPsj3g+yH3KtEM
GsJMJ7sZHL+9K2BXIK0kwGOYUa4wf3Nqg/E4RrH5MFV4WUVDHiehpGHIUuVGV5S+8TxE4Tjv6iBa
svDGVfcX3RL1B46HQfi7oAdYGP+aLbJWwzpIWp+oNPTRGi4gNMr9kNv0tXttkmgnQ7uIpRggR5XS
P2tb/HmDvrgeZLBIhRrD5xBei89jGSPIqF1S6SwOo8S7mNS3m3l2JJ7KXyXq5WGCetodg8ztc6x7
BaiFyVrTyqFJAXTnuyq8dpYlZ4IIWe43d/Dz8mv5uHI+Y2YLJ5iYyrL5YVvlX++v+1EpQ8f1I1X4
nsdLBZcXQa7iJrqLKso8PozcCpANRg3ZEKRXzUm4ToX5YlKXtAb/Qj2TIwYzxAx0CjD4jzDyoBIB
Umv/MPGUuJ2upvLf8rJk5y9l60THgrIdipjbXhh0jUJwEL1bRQ26zdp6xxWxe5V33icAIoC+9tA6
XPn6NWSwyeJ/PD+FMk0X8F9UUPD0WxFYoAeROAKir1hcjEuFQAsNa6ykU2y3Krc0eRnnMQn1D57I
ZQ9On0C93vX1BJnjBUAHEdRanfdJlzu51l97AV5ow03DfI7zVDjKIxE7G6q1EUCT1aN8J14NHLbu
0X7reZCNuOyPdsPq6yKI00G4S7PbJ2x8SlBbFjooSTaES4+og+CafhnRh/6L4OLAn7TnfsyEywGB
24YcA+W2FXb5XbyUHat6Guw5U/9rNVksT8hab1zI4vwVUo/l9wDxEOUJobqUYTdxgX60QU4xbhzs
bGPDYGjwpirtQJttXn/S3hyW2ZdagB301v8sPoH4UOza1kKnVFumeGV58rhnupcsDyWgliW9AUyw
r6GScjZ1ZxQujQDfSXZGAQFRGNXHZNlCVgwrzcLoxOre4okEazCsW92VXdoROYDJwGqkypJnTg5q
UpS9U+D4rCFq2Hx4o4yQLc1n2IwBnoAW6ENYPltSj3U/TmfZtZq3trvA0hkSlpeG5hvZM3fH6iva
onJ9qmjbUz0puQ86Ffn5+cDGXbXKm8xQeIR7kCNkN+HS+/Hv3LfkJWYgvSs/w4WxmDAm4QLx/jr5
cwvEjZxwYTlBNKbrBZ9vykKd5REOhOLgaW+sHpL9trnWOL+6WoemSlAe4rQ2HvxtHx/DNH4RJBMz
QsYogdIQvingKpxdnMspIedQ3zJBR4Y2mQMuJJHtlr+vQlDV5UHArr9W+2ucFDJVOEwxnL2btd7U
wdkKqeCPR6n9Zxn2ezuZoj7JQqLreW6g5f74VZE6kpmmnijFCCXgWGgeNsmm6/ztvQQSQW2xLK2M
GfVYdQTfl3//3LcU5JP2sFuI9urtr36qSTU0VnORWH6lynR+jHfH0bnJRCiM2az+scXUKkMYAWr5
4AKlSZJnbJShvWYfiLxMGbBo5+HiykajOwJbqB3NNN7eBMJJNkeMa1Myxclm3VH/ml7WhSkv/IL1
uACt+8wTwo917KAl0/N+bjrQ6udxJMqvAaS5JPtuClLJV6zfysZUcr7HY3BY7xX699p9tzrO31z4
8EflysKI9CJ4hJGKNwLiY0uvMoN2XoDcJZ0J1d6VQvnt1p4LXDzPSFNgkR6TU8qcJDLrvnC7caYG
R/bDwWPhWOA7HiZvijJSqQ+HjmUXklXsSc0qaWERKIA/vq6c4qXm/PGlhndZfYnZjzuxTUgGGuyD
yVhse3ZJe798gyBJhVsihVG2AfaCVRNu1tk+87DvLryE9hQ61+Wr268nqQ111FmnQ0/Smjzyjw5g
e7PsuCnAmOAMCzrUxpXLXNblQuWOHIWd0JZY8VZlhJ4ZoLCcTnbnr32SIJPR8zjjJpI2kA5DgX2z
7B4U/JASUTFyPYmJm5mCAGdMHQtFKMzM20pi4RsVoCmEiXW7bPDyoIi0+BBF2pN80FldSqyEx5mG
hPPBaMGsMgP/XoPjMnXyvsChSL6E+kNsCv2KQJxQe3CuJAy0SwbVgM3vltA1avatNcg8h8yAI6cc
dPay7iDCZbhNDB5EwuPxF5iiA31Mmx7EXAIsitlUUToUb1106Slvsk64wlKA81ZXf7zx/Y6pG+5M
xMpA3QkTe3DjLs8/mdw2rRjb+/4O+O3PkNE0yJPFg+JFJE+eXzSpGLRMCmSETWjgkEzYCUE4mGk6
QAkTNxcSiHvPO866qggAEjZ0dfqqlgtyqeX68RyIO9RG4ilSEydcqedHBpVaYVXcGKLO469P9CTT
Ows+jra/D6eKB+NclfCVFtcojR/csMxaAadrvCERZsMneQAajxehIMAC+CMGQwPpLlMwPNWTkVd+
zHGIwey2gK0pECZZSJWStoqxmveud27+zbaP/augivrl3X0ldZc4iF13LafyV7SzWXIr4TIJxJux
KyNpw3yLXMmg6ES7mgVIEfLnBkh2y4vRkzRbkqEhypr+/eKxW4p02poIyPEk7dFDfgcKQlhnXkPt
DbWFJHOKjRAg1k11Ypzhatm/hzmSIs7ZddxlVmjXxihzQl4lI8fwFFkNCZk00yU14AJZ6OTugvOE
0kZhIc6E6/ETX8bs8ug02LtpX+z0tssOQ93Em8W0+pdHBv9D0VoW9itgcqIRfUJzMuSKRveNuwvQ
g96IW9dYnzRacfc3CcfU4pbj/WWiETc5UfhchBJWaO2ocX5rAitOJnxBsIj0y+h8VTOO65mVyj2K
rmy4KBhrW9l28EDn+qFzKYBgu4udYHsY+9N+e9osKeZ6rBffDRcV9U+U41Ck493D5eO/DKxuieoY
imWwJHG+FJqk7rr3mbVOdDs9+F+4cvkzjDHD28lLdzMGoIrnr/8nslDtIZNCxBuIEaI5DUDtTUGe
xBzTzMpsUFOSrjQ1Ox7Lj8UokivCTEc1S9GwpbYldJT0/ajCAhJ3FYZXqoiGyw6WKDVj+BbdMQVI
h2nbET7ej43edIjq331GEeO/QRAG2OgkHnSkJgDKfVum7uxzYjW1/mowISjCB4srIbg9/q4HM06h
YViPPNTTvODS3jNZyNKP16n5I/EuZsk7iBMdsDHVcrB+1XISJ1AVUkfqO+6eCMlBAWJsU0Esp5kB
dk/h/81JPVzaj9OWT3c8zqnY6KaFgiDpi2oDt4BNhjTcyOHtqx63hlIZc/N49Z/R+F64+lCJ2MMt
cs2txqx4I1tXmFGfcj/mvRkVMOZI2D1StZz/Es7GyoQeQz+PnT71JUTxmwuOckU3yKgDmxo29FoL
THckX9txJtb3O+UOEZ182lK85WP2ZDh+vVvLqaq/Vm7whSu9Jz3Q1OH2ue5aHQTfxOP2femsWjHP
MSvx5+P3+LFvgtXuzfBYEUD5AXVqINfRVMnCD0IC4FM+JqRXOfdTwoyauxZyb/P6Zy43H1oE0e+r
+An8VDcefZznUgn6nPUp2IjpkhwxEUrtQqhFLibR2k2iM6GpBFI9MEB0XUxVJjVab6a4Y3TujU04
OUboF30n2Gw/4Rrp4wdiqvjf66gs0KmS0Jlb5GXW76W9oR8ZsE1eif7wY4R90Dqoie+VDqsWm+Ia
Hy0CZHJzwJoe6uT5OrVSlADNrQVbESjBcS+Brp5OzD3D0aao61P7zBRSK8AZFYU9jAAB8Q/cAkH6
QwMwWVe6iZImCKlrHZ3PCPENXGPjr2WSWg9L7+5cqmPu1CpqZCrsVphKSyEjlrlQQzs7Wcs8WG0s
A24pyd7oJMxaaYf/bZfwt0AovGUPFlJkvuy6ZBQU1I/NB92UTndYUkZHx6nkGJApB77yMN7lBBPP
nIg3MSjtXCR37+o6ID6ERdOIzzcn13GvWPu4E18s5PKKdZ9o6Yyny7/CbBMOR9FS1VGAuSehM4ZY
1aKbvvSHBXhnR0g0O6XXV7eQgW+L7U6X9W/lHyb6sl52+tEaWzpV6WkhBj3l7p9dtp8USEDvkZU4
Sm/tPp7kSiyXC/kWSpcNtYB7+C5L0MCFTBO4b4f3/1ZvVYb/sxPboxk+/dvue6j/mF2YQa95BSFv
qoFrASW7xaXsYAYiKjA0DGOdWle9vujI7ZIE1LWgd26e33gnndxoFNkshyuBORg26mtDO92Gs2Co
VVtocWvDQ4GyVZ8CnTKuyIRJpejvwmgkb7KOBsAfrESCR9rKpnx/YGFJ/KOJtvouIro/jeuaMIVD
rb5gq/YmHfNd5PRPCa74grf2zXvqsoCL+hxGt2Xn9aZIA5TnF1+kCHemjMfSUXRiMXZEFvDO5/Iy
DhxYAMlt9Z4glCTcaeyhIvVBEiU2e6zkh2OGFzTM8U+GPXpyzUPOeTp6OazNc/LFrHbt0eR3WzKq
J85c1nYdygohfFj7HSyieWNSye/7B8tnOIeWGDpkZU9jeSNgvR9UBK0GT6l+ZIEeWA5gXELz65Ev
pHqRzwy5gei2rmWVXRdLrqSaII12ToW+zFAT6g5V33nazTyDDW6gXSRJG53SNQRlWsUwOYdYO7KK
Z4d38BeX1UrhwYcbX9lB58q4xZ+ECQQt9LDibUnkU+WSJRRKtvBWYkrwJuv9kKrj8CR2LsxCmy5Z
rUvOlOfYlJak2u/I2gIDC/J70s67GA+sicL+eZAY9eNNjGr1oWGYxcMbnFT64uelkLEbssiWfxes
xzMTfk3f/SofRghjaHED9tuOSBYYz2ccbTh5+0gjrUV2hywNfPRNchNnMttP1qEDfna87VfHAWHV
JzXBcLlo+8snONuT/Q/kGBmmvKg90AfR1MX8cGpQ2W1F08+/6APTRWQMzViu7AVcgC/VHw1Ao8sq
nHNRlm3vLxpDrcIAo4JzyDf1GNL7B4kdRSKSVMpAfr+1hc3zx7wRFoXGeWIhlbg9uM4/4GXYkQgw
YnGn+Tkjl/OX3r3rNHk3B0OslyvUVwpMdYR3gM7C6m4rletgS2KzORlSaSIxfwLHf1uYQZ8Ye2Cd
j9lKAk77wP/MUNcgWAg9XvMDSNDyjsB+y0eTyTkn44K0i/vtpM8Lt7zst6Gr9zbGJfXR0564IZj3
1l/uN3HU0vXIV8KUgjjeVYyx4i8R75WDEXOGmIC51aGmlTHybH6TuyMjQV2RbkN5tWVyoko4+KKJ
fkzy1kQc7UFn4UD+dpzne0Vf4bslorYYlCMTsvu/4nDbODY0Sf/Nbpm19Fi7S4Rlkm0xQSTdjhH6
v1mka/c5jSQvvwz5TFioL+EHx5Cv+Fs2D4VWo0XWVceirrDATLuoCkOhkN7SoZsbvVXWw2OkX4it
IxLt/bJzZ6Y8E89I7obE/D4EzEUbVhZ9AcfNCZJN91VPp0tEMhO9go+G404t8cJI1GGUdAVAZleV
CTvBfR6h3Wd5fSeiF4vjksMpJVK/PlpU3kNdBcJITLKyWuOc/PMNiCF+yKoqZf5/OObwj7wYbN9b
ARd+4T3TQNbGhhzWjtJ2DBI2ru60OEoiUzApIOxkxjDXAR1IjwJmmZ7GCJjamTO9gpn0/UHhbCBO
rYJwexj3bU5ODJ6lUQ3MHOBRGCwlrN74rnDpFXtd67MDv4ddQpAqT/k88/5xYiTJB7tFod4IguYt
mzFgzHb2EIHsqsS2dO3921ghwbT8HAmdM5dOzCRG1FhwKOGD+Dpo8T91NqtH7set4X0+o2WcJgVO
zAC1zT9OVr9wQosF9uAiyxwtZT/TnZTXpIElNqHAznaWiPGM5TijV1oL99YDOeRRhwxkiSjuZoGP
raQ9TScKt99J+3efeYqxlG92adlLgCSTIvY/ChFj/lQ8gIx1nlbkuj8y/KVEIUNNxKhALw2ErQHG
69beKnyRraZK4A9JN/Im5NycObb/8JqMFeADMi0UfvCg6MIzjdPOQ/rip4RTPdVWzOETV7127v9W
l/hkc3tZLX+Igj4Fc/Cmknk4VoGgJmB01Y4w7hudx2tdoVOq2zUJE1hf0K8vfGKQLUistVOaIBRr
sJU1YIM68bAulfyrPPMgHQk7XB+9ZU485cWLQNWBTmKc82uulc/wZyh7ELDgiHBMUh9M9QFmnaDn
ptGm/UYGNc7b5wMTZJ/inTYONJ33LHs/PG8moGmcDm7rcL5cRPS7LalhB93ceylE1ZpIERmA2+od
ESXhxwUnCemeejs10f6/grMWqgAoQ0oo3AWqH0N7T9VG6spnRrbEkGDHgCygxFKS9qhCPuwjTw8G
E8dTyYaiQd1UYx9BAYSSggihl9fGJmVeflBXSsSz3yRwYeNiLh/0iBWdYXjKL6UMRngznCaL1tql
uT5BwDlflzXibxrzzquFETojcGAHv7mQ8IVADfNxVKhVxHO5ieGex+3KoOv/dgiO+xxL6LGjjFlJ
9x7GeJv4mrjMRkzrvtLkbjDNtvdFh7dPEAyU3F2LIHSHdl1hgIrxzKhtaJvtsPMzYx5GViVfucVQ
JwpVsYOmzNu8RTmiaADJa4eLRwcoag4SMaX9tXYERsIKPiRd+/uDrHhatW1bWQzfTJDr61SoOqhk
T1eIKcCz9eqkNujwyyG/dQaYXg+BFEKgW6Bg7y8zLvGI4y69gV0vmv30A2RCGpW81GM62W4QtIst
HRvj2iPDKbUdkDnpcGalKroW4UBbpaYJgXnpQJzYwn0HfIdfYJbnwCHnP6hsGOnhfF9LkMk2lVKT
HEHlYDBT+JupH0k2j3BJilghzXizipLApd1OYO+bFFkFSP/41kitDxqdjilewRdKU3l7XzkZJChQ
nMCNxUmViQJurYOtQ754ovsnBqC5wii5ak4Qa+l8q+MJGPJXrcSMXpdTvAmXBTnC2XD/atADFKwe
RURMuo5GV8YrkoiJPmZhjGuSLxWYFU7mXUXUzrNyJU6/jdG4w/aNkJEWNd2pZfb4wttunH8ObTHL
wCfMcHJlr90qZTcbWFwPe151WDAl3bq+/negklNotBtbJFpK4n2mJxKlndviSh2KOOC+asH8Eulg
220JT5oAZPbOCUrsF4eyTRj1aMifhBhagaXynEboLXREiprwWIxZR4wgekxFwhhIVlHnRdOMEOx/
gYvrtqkAMhO0hF1SXLQUqaWlc+7O2vod+FKaHM8PAd68GRa0sSU72zEccjTCfWun6RjEY88uNFFw
1Pk/4T/OzvNMtexDkpx/+K7oRR14lEZFw32JCSS9w3GNTCPf47DB2eZKzWqns083ROupTtLQ58F0
XOvePt7GVucSm9BKlOuTCevpAQoD+6naUeSQGhX2LtlJr2DuSCjg+8SvnwHweKXgHBVUd1xk454V
OMVl2Zs278tvQ2zePfM/dqLXjg0I1k/d9Ndh7MruJDZ/6LJ2MSF5ziTiR5jRUmyB4K3KnG6W3XVo
OY4Youa3tLcigRCBXvygaTD/t8iib4LLomj4FWNfIZeM9iyRWdFVJjXFqpUoCVlvW9gbL2m8cOZi
vARuXqOs5+3m6m+WujPMcgM/AnOkCX0NTTQppIXA10F9lDD1CVQXADOrF+aaYQIog9XuTztYb580
9/uvfuDB8Gog6ImDPHpmKhRyI+mT1L5LVWuqTsXwxwsn12pp08a6K+r7uyuBXCP+25E0T8rdNWN0
/np8P68zMvQlZHy44ZAbuq/tkqZ4h6UMYeN6LZX33lxphzpMx9o4lqolltS7DE2/QWZV5R5yYIVY
DENH+V7LNp1XUg3EEVnuryzgzuzdx/DGhsp+FoYVVUz+dsLBP7ppjZx8fhRpP9rNQ8wgfMbF5szc
q0/Ihgizqzl7zdahbjA7Frii066/OXZReRs/aR73b6KNERUZm6jlq4GOjz2HWtJurPtOCdsXI32u
I8mMkQYLTshk8Ye8G7mlyG6LSnPHHseKwTpr3x6kby68fsHyoEEFsJ9osdCMxRZlziprCVsuhSYo
5V72MyEZ7RqJHq4amxk6SX33IzLWRiDsnTrn+dMmYTfAtgSRlffETOzbK2q3jU6ywof8OFdpkT+W
DgwkDFDZLuONxE4E1yA//lmPFOiao7Qo2JZysIecbP2Ey6LZ3rFaU6Gbzo52PCz9DX2D9tZSUNL8
U2VVmuabul0Xeb85FOOqlU464wDm6hQrTkRWUjasWuYqDyqDvdcKL29a0u71h2aG5iGO0WSmpyJR
pvrSx7xGDGNyIQNXNQ7siVnCJOWlWTAgvWJP8J122fwSEbERrHGjM6Ob/a5MJ1ecvcD9exQvkuTx
Hpmhqw4Dn4aC36hdQPhfxNJeG+qv2+ZCaClJiKi0ohwlzx5EpO2nPZGfCQzvUJkqyUNVlBRkKiIX
aNnzIvrDPolm7HdYrcs7W/De2rzY3/ypX3lKQUnijZjGs2bns7rUnrxOYZr8szeNNkoJ5n+I/ApE
RFxYwhVbueCYveh+JpVopP3RLz/MEHd+Q/5S8AIPZraDWxiOnBUtBmVAo3OsrFEZycc3McJ9939E
3jfKGc5w+fbUNUaMKdiOqd1R5yEy0iTD9rXudKNLDOAR7VrKPmp6wJY68X4BLRJR0szkJinLzvJE
0szXPZY8U4ya5DaSkYbGPTeKFKJg4RXaVNVQb44GkmT+0PXqJIjf8+VyXVO2fNXmPSpFzP7/+xZ0
H3m7QCV1khSNDn8Te2b+KVSLo2MQnFchE1UIRQ8bpnIHbBHUy8zDcj+9j0xeaZX2OrHQ2FiXCW2B
NCFwJpwfWgfKqss9ocNt3IhVkbLzy+c475kI8o5M+nOJ2t+W5pSbdejRhNbcTgzLEMt8QsCtK6qp
eaGdtgsW/WeYZ8oo2Qjqdb0mSlgX/aXn2EEQ5GQ1nRpvyFh+u6LHnBjej4zXaA6PWG5Kr5AG75GP
5eeabOwWIhgW8E+bjX02aL9kcsWOtS8XHmCrcBH+zzWBuTvmneBo0AlH57MELq/MhZgJTAvszTwQ
e3pUvP4nfuTd9Dfr7a5c8Xv2tYJq/+3NN9HD+Zdillf0EDfF3ib6duOPgu2NLllSFoOYG/90+UCy
TyHtPS+eXldllXvCzeUvD0l6AxpB8LqwTlA1hs8SRfwa+zxhmtZyEtPduaaMYupF7NyrkpQaogsC
P9KDQUNMYKh5arVgFPU8Binas0/dQeG2ZEipFvRugRoV/e2EemB1ptzNvcRRylrtF3H/XZhxgi1I
54IWeHsxNbBXjhyDfFi9unfOLndjTrQjt9BSn1al3pm0wQjNsIffU9Jtf/3fgmzZXmrNicBgilK5
WfD5pbOuq3+qao4R0CelIrjXBy0A0ajS3KAgzrTIizBEbEVP08E6D0ELooERpK6SwwMYCH6A+dJO
i6/f54EfHuEPvc7mzktFWwhyuzCBYNyebTOyRJVzEYPQpRuMIUbiKWH3T2ds9uzmCaI8d39EBBqW
gMNhoAsSxplc6u98/wTAVeKdxu7we3ABa8Flv9Yk+52UZyyvewatvwgctIPG/11hw1Df3GsXG7RQ
jpFHn2OHSUzkPWRCapJ4ARClsm5XYDHrXo00YH/WFEVygjBrwGIHJKsIG5xtfTdR8iTa/lQg18Ta
b1vPvzQsNw/sCi2EICVa2hm05kB+jA44GaiDy0xCEpKgVqUWx6cR1NjreYqxqcnSqTC8DeG2hlRG
5TQjIqXqdvIspiyle2oeZMupPCIQZs80iVZpvtio+yvSDfsWejrQJSQrOI2sl74Ld6YGAeSesoOa
GsrfSmBMLzpf0WUwzgOjdeowXOiHr18dC3e84nOS5+DPL6hy8saEYfa+YfD4+3C6dm7ylbuidYbr
KobbZMgC2+1pkDil/CFvOCPQaPQDHkf7eERQ3HurKyHpHkyWUiFrz91V9Qa2RdcT3UgLqHwpQMke
cDR9XTz8WY2bAL8e+AkK941HD+r5taUuvDgG1LDVFKWuB+09yTJvMxi4G83bYVm32wwFCYZ0pocH
3bsuHMzGeF4ekrkc5BlU/YeIarQuUoxWge9g2Ueuw2XXqplcvqBQ3JUP/KPHFa9J9U+RsQpoIXld
EKjN5TAoAbFxTjXz2a9w01zJfqZSChAiH9h3TPpqWrm8xxvPa94tatETLURS27hk57ZPLBDwdrtq
T14WU6xPWNpo4jCi7u96DFCQLTNt7Dogphu4cqeN1J7EU/748GmIuWx/Ol2XG+7l57jlXjoeEWy7
uycenPq2TOIq0X00MVbo6RJ0tPYgO8XSJlJ82hwPBohOh8qpqKjZbw0tWsctWpm1Mab9HciuWeks
ciD9FWOdgCNjXUPH3OuUdpI3jvgpUPg3G+PDUKueibVxa2apwTgjmpxKJYpwtkV3pU3F5GRFgW4l
QysYLYGC+SHXnHdD8ZJXfl+tyVa/MdtNxX0LmUWNaUB2mal83nP7Bdboi37I4qGNhEWCfzleiSO9
KFyhV3pefTmaSQ0ZBfA2b8yK3lr+s+ALZhUVVi1Ai8IxSzn5IxLUM1Zyiz9PL6YcVw6Qpvz2n+k2
s2bW/w4U84gMl2GLGdGYFJb/1PIRHQGBj3hA0BiQ1jBc2RkCTZyyspEJcvd28DoJA3Y6L0po6j35
6EDYcug4CCU8a+EKEqTjPNYYEv9WUEFdSq7LtkQrvrPFbmRp8/Aujz4M2b5uRp7TRjNfaTC0f0O+
Ff9xvFAThTebnDFOIhCeeYKUEzArtmjsPfr+uTjCnEIRqBQw4TjqN2A5lxFOIcL2y8HpFaPkeNbg
BNHkB3yecVMz6cyiyyHpLjf5RJexAaUIrcdMZX/o5t9TdkW2xWy72yFssTcr9wIp8Z6S2aOiN1Rr
PeP2xYXn9h/pNAqAY2+WH3PxciZXOe7LL5fhEJqLh2inMdHcvFbeYyC2bGiPBbinMHjIonulD73n
M/nH6SuPbbdSzs793HEYwQckw+CLr+Xa1hK/DCWBe5c8EHi5RaFUGcJUYZ3JV/Qoijx0IolWOxqe
827xUsDTwVSQcC7O51juZ1UxiRPr6/TfgXbQoRJDmBgq+jOZqf18NcDPx7Odl5ZDcVm2+YdHj8/n
puI4Z94v0AFHgpGi147RkJS3bV5bevmtJSmlfNW9fowTeHRSo+6ixFAi2E0bafIVW1cWQo9X7jfG
wmT94wO97GhT74kXWOe4sk3zdASLl6YrDBGMY+uAglI6ENTgnaWNOCFBjsNbGgq6O+aOw8cecjPc
aRKkueY4mjCX0gW/RrI8tqRRZfe3AA/j3oE+tDyki5LGB6qRpkKwShPyFmJy3zRkS40EMyDqeeMy
Wf7hzP2pKCSYK9ojw01Ko/oM2rzGSDbusKnkXYEXHIABNa5W8hh6s4vIuyHA+Ca8kqNe0gG+UjXg
rnyyOZiBBOBE1SiCFJAoaX0R0hmZFc9m6jBTzRdJ6k/BOdkX5glZNrez7JtqSpdHIHGEHacXmmA3
ehYTUqXKIr26Lq4d3wV1Pr6JyVy7B0PCw1hoRkzspVvYwDoGgrr3JzVk4fii255XALZ+WOFSl3B/
hesGW8w5pYBRohvTzeOnHlogpbVnm0kBv9ecC2maL8HimfnujxIrk/hjDyAx31wmXyzXc3iUXEEW
m98NM7oIHT9II0HB9JRMDHlisN5DXHyRe3zEx3yQgRLh30Y56/t8RydHqTk3UOHWpM6hsh84nn1n
Q2umw1bzEO+5Ka6akFTWqhqNjuJwmcEJR1esvhmkSVAjVMMZ6lmuFPgySuTV6eSaDASWaeNp5GYy
v6PKf3gGh7AC2aCaWJkian9qLAzItZ/f0T+/mfTTZbU0lQ/cAlJS79K7VWhjYml0gB3rthAATzSG
Ai8t64K6NmM2fcHffV/pu8JkmeexNVToVgbMd0NChCga+KugQJnhnQTlOHlI5nFHwTrWuT+W0fyq
x/mmbsXWO7N7eWJL8ARJLE8UbtBeyivfNl2XEbdHOnxUN9g17aloFngugd3Qy22vUqR1HtN5slQs
7wFumSO/9TgF+nzHUqGqnOm0CZiNNobQsgcKExBLZrvE3l0j17dCPw+ETpWErWPyevbwIVftq+mP
Sersftl0f6PUaTxFikujekm8enfCn2VwRLx0LOpNjDXhNDVEYo1KzMIKG+gZO5GFi6p+ZsiA/LR4
bDv90BT0+G1h2RE0GhCVrJ/NVp8ZvdxmRMl5Ie22zX9xn/eKo8MaYFNciDZjNVa+lHoAUl4eYYn6
xw5pMhQV94TLnPNBj0xvbBqY3dA45HvfzkGdaMEiXc4L1ED4K568xCKBDv0R2BuZMUXNHLksnSqg
h/NXOQQyuG5vTv5RlJPWAKYenGT5hEz7AXX5mRyOPknlynufSeBGHHW31alWy+XX7GphUKUz7hZ0
sDP1pPKr2u/fcOWGbi5Fog70vyz63tPBDOTeBJEoZpd5jlmkdKIx5UZ6BBPaeskwELRa9SRgXexL
0gUHEyV7hqZuqz2+vUmK/+TEUGV70slfwAgScwZWzHQP/y6kxtEMvRHjl9avlxFgYuRUPMV/GhF7
kQ2+t6WtONlKG2LxB0Mtaa/TatTZLie6gX5uNpph8rgNNmXJwZupBoLKJCZcxRNGQE3Ju8SdZT81
cf/MTgvzrE9Of9Bd/em+16nCF2pF2XoYh0URfaXPF2gEJ08McI6pk+X9ECy9Q0ZpjOjKDvu4Lq2c
CMZgYcinnLx4tEqvTfr0Prd8eT4/T+4k41isbfRxRQ4zm+SJ2P5mjl2lfqiuMwic62vfr+J4yhI2
zLWUssbe8AtzKpJzLEpS9MWFFCXcVyUNzqc8OvxSnxbdH7FGN5VJa7eJ7xOtTRfz5ca9GuK/y6QR
M/dPPGPDVTaS3MGtAtraZtFepPYzRiMUSBehKT/dQ6BJRrYkFcqmGu+ew/dh7O85/N10u0YwHc2d
j7RNCsxzgMgNVoWR/zuSCe2vhePi3MQwC4FWg/ZpQbLMt5yA4fqgw7TMkbK/b1zA3BXSRcbq1EA0
t+bDuxu+vpG8ph13J94BdnXrx5JOuEGefE2G2MXpJbxRehqOZAb5aAVLL4SWS4lE5Lgjtz5wQ7EY
UAy1Yj5DK1YVU3DgtuuYgPMrxqxuoxxKbX8odwUFUoZFc34znKYVqCITAvqm89OB0kEfCZl3Xa1Z
cXHfvvTeqQg5a0XEsI5b/yAd2rHafrNroDrv/NXKAfOIaBFFY66ARAQ2O02gRLIJ8mEJ0qHeNiPe
y6J4/9gMhDqfNXYuHtEYMz9iJ19Thl9OeJhK8t3wVLUHkjV1xnWlyQQaiV6Up/X3F4Ef2iMmMTwa
LOchllwjpiAwgJUBJCrVNyVmdCtq0HVY7NUuO1/TCuJn5RhzsDu5zEM01R8nSzzNQQRgbgrbDrMp
BTdX/IQqIeXmLNxDaWAXENrrjaIiohZcf/W4TRpU7xDJ62PWgqxioEv65u/b9QltWG414W/8e1PH
pzaf6QTb9+c2vdhBUYyAlLPlNvr9/WI6J7kf6WNDX4tbH49Gk9M6aO5hqMDMrMXOD8E5DJrM4pao
VZMljJPlzXXlfFtDl+YqISztOCIGUQT1IhQmy7K5/4WLIKfojJzoGNXJWozNNf0u2ja8FUHUfsi8
OmgOYs+9RogbxJNM7LNXEo1vyHHGLfVpS9PsSZb+EHPx07VBwn/Vq+GDyZ1iNxhLHHCJIQpr88Fe
OoFffFvBVHmgFoED2ZcxDKOvRncFe6Y0lD8jueGkN0XWMbQWVg7zUG53j1GZmmTK5lPnTqesoo/c
goq0riUqB1yvnhLx1ro6gFhjhIMs0ftDjGjOyBkHlowMgVa1gCJLHgXEIwP/sQwj1L1jTJNveGAk
KiBivMUevAAeYiEdx0HIA8loY2/bh5xc5kfKhSlKnYYeReE+tYRYiFnZLVAhe9sxDNy2HKM5zjsd
FF6bR7ZxEzpm05SRZeCO8F9i2GtdX8z0Mnvv2WPZfiOC44XRONwQC3qTFaNn+imEi6n2Tfa6/oQn
AgQof8PUJ69yGIMIKzuKFzcmWLPr/0JwXgI7gQAoz0//d59eQicUhBTH1nWBVTLdGdgvLecUFBZl
P59YS5EC9vIVtfaKYILWj1FPcKYcr6ktke2iAIc3HRuDKW9aE29n5IYSp0Z9QTnbR/JPLYJa8XEO
oiJERM8zLqhoalNg1WiV/oNrh1YNezYSH3p7HFM5agvu8x9ORlfnC/1zXU3KzHDs7QkdV0iFY2xL
YQh9PldAPRfH0CZFroOwXBSpyBQJcCagQ5yPHpP0QeUaEo9jPFA8emc/VEx3qkKVxHpuppsb3YQ2
egr2jmx7dB5QniMgkKntYWaT0OdLt133KXM63LdjcQt2FHiw4cefJxGgKHyHjdC8z2AFCq+YyQPu
baP/DUS9ZlL4/t+xQpO47a+nBpsF/zwzOu9oJA+y6x25cDOY3F0vTXQlLKjtpXINdcOwrlHys8zt
FuGFUKl4JJ1YR12eqbFaYNpQ8THm5iMpIeGXvu0accz14TS5tPygGKC0TMrkdSwOo+w33AP+XgY2
5eFczqtd0GkOWVdtSTLZGx5Z/d0K2cCevE1oC5icigc1OngY5kpY27cqD8YsaK4i+KERnb3ZMfxG
1VrSLObxbDNHVcfwDaOYVPyHIYvTO3vti9naZ1+ePHwYF6NcVfNwEowBEp7jl+B98YP8ofq9UJzo
nnyQiigP1LWarkLVFZ8jNV2+hpvwSWVCT9WwiUwaBGPptt67jjwPoPhqZLDg1pwwN3XSXAGnXb3I
5gFfvDhTy3pSesuhU0kHzmZ4rnC/emLDruQYCXh4mdDGhEjoWduoWG7NdZ1mIlNPJtL9oVOZ3SBC
HHkHBGnLN1kPmrw9a4rorD8ngI7gefOu7Joulz3wiQG3CQysPKBp7AwME6VAB36Atke8dKqvAEJn
5eSzjstKrbhOQl1Mq+fCiYl0kaevkYGb7RGCzdRXXcp8xWGHRfn///iuI1utnIAq3zGpHCIgKLGr
yjIvlbAnAQCIoNSEpwveMQwxOpzd8LnimulfOlAclsxM2McYShdGVy58u5haEunw22I39gVlBlV+
5v4HpEuwoYEIvRKa1eMPkxXsSbjODESB3chVZP1aDBpbG62cDWR61lyw3ELvYHG90QeSry7hHr0t
3UhFUIQR/BPVirRrVhOrUp2i99qxCes8pEL6DFNtzhuVwZvB3aHTGM1uVxRzgFxCRtLAcJovIAve
hh0aLJiopyZUvMuniWxY/2plG3EzriYMpOOPSieRwg3hajdidGLnV1s3fsnnMsjClI9iGlsSaLlQ
siYBocJVA8mQJnV31boAR1+HfvVuuWTq+DHXU278fLX3N+M4PfOghR9tjnBBD61gmsPZ3Mwty/qZ
5O2qltbrhb6ODV5PDngYmnXAsHESb1kz/dEhCH+hkCreOARSRW/egHV2lKOqDHbNlWgsK9qnnsyg
v4VWzsyRylSzPhltajfUFjhq1HHhVaduvQV/qfVERIGD8SQ0JuWs6AQMvnT2gICBs2QxNXttpp0u
UlSo59Lxcp6v7+K3s12Pli6BVE+TodPFCnZBFy335iBFx64vBNnTtRLhvsZSxrt3HUFBxf/+l/J+
ie3D1AOGHUHlNUIwZMYRSCMFPC2K1S/WuMDeY+tx+Jx5fOL8BquL4tyunDzhg0E3l7xBNZNYonQu
brtdFUxzKaW+8bHNKPo9g0l+SU7nLjTjukb5sHb+CKI0xHbOlspPUB95kEo5C1RpK+Fu++q37kZW
tk67iTETMk9cDi3rN9fZTBllMwxuM4OeWLz1GkVgyJsjOKtlrMaqLVIaLHdYF+XdOkufrPiBHzgV
81qeNdHVuAMS7HcMFks+oKmRKQiuVPTBuJPKOuwdSZ8V04yUDv7M4DartJIVCVtV78dElSL46jPl
c6bleq/V6cyCg1LVgijwDeN/7gMmtIDNm3ouk0EF8LzeTdmWU0S0wm4x9F7lbKU0E57MSk7rpdl2
fbtPQkHwsU1bKIyBt8ProbpWyYm7iN/mqy/2b3mYZL4nvnzyytp4KBsUqUbTn8hHCYRfOlwcyMFB
9IKUMktthWcr/1yGjdt3QRteBknal8dHkzAyZ7643GuQc2VhF4u/5odehLROUe/6h26aaoa0ATi5
oJY8JDPZzLVkuLrPhj9BPaIt4BsDZm6HiltWY0IY4Fmdc32VScyptt7DxSeT5WJzuiycHyRcPp1o
eg70pjT8CGMiInrgajJC5+8Ynu1qe3lehjXD1ZodN3cNo1OYO0NywVAJgijN/SEGq4zVd4Kz4HJZ
ooitSop4s5jk1ru04kYFmINxWzFWN2FjQuB6++tPpq0KKEpYbejp7ek13g7m8wZLfRg2r19uOWbo
Cq8svxv3b4u2vEQw1LtCf8jRx6Hjyf+vKrWQefN9DLwUKtvhFKZ++Bqm9LJwjxgrHdZpYsUc1Ued
iOO2NS9dh+LBJV6bXdkpzzxGznlInVyA1n9lG/cTbgqhCGX9oCpMMyGZoqWL/EsdN+Dz9qQvRk+8
xBv6E92lfDIMCaV0Wqf0IhqPSsLeJDOv5m/wRGwzwMZDOpmsUYUnXZpx1Whbc30tXb1iM5KmGMmq
R1FC008cSv086dj4q3CLbi5lxp9l96dwdAajgQLXDVfYty821UIaE4WvcB3pYnkXcsUKwYWS7hRr
29VJD+wiebeA93wtAS1MBTxjS6YeSwYJt5lV73RCqiWXZ86lio5ESGSHuQvETeoPEI5JcJLb8jNu
00ADSBt0oux26ZGZn1jK+mgx96Fqb6Ep9J35Bx25R1dgB0NxrnwYle2Pmv0Nke5QonADtKm6vS62
ruU2kt7wxQGJszzd3+Lk0atRsS5G5HwCmIDyjtg6CvrzT7sxdl1vfaCfBa1jt8FNybbYiROdQhVN
PsNKeDJcERFnnxWtbxa23xW+Pg3zAuAzsXclD9hOjK/+tdzlt7i4Im5VLd9J4B7HI6UVwe18ctB/
uflDlFTxfw8odbXmbupc/wng0DSvSllkv12OywiyHUkxEwGBLAGROR5Y6x6hKyoP61Y8MZI0L58S
QDSfQxqShuJ8zVmrXCHK2EpV5oN/lvrz26d7VUcztbeN4BtiLp5owZ+OFapIBHdmZMu1ITvy571P
x3yxTAb/ozz8BUJF4p53HGdn3JA4Vtt2Gon1Lgn6trtchNITQ14mQMTFnNmBBDW0TTtBVWnGNhtq
zktyWAdZcVynGiiKZtjZ8C3Xt2F7Po9nNgLQZI/hCGheuF4G1/TTIDcn8GthFSsaqXlP9BfqlIG6
MXgZlHIsMqb1A7/VQQ7mDQl5jVT1NaI3x06PFzDT/lL8vbf84ctwszUXVxsupHXSOgDDRbnoa8bs
1hHfwdMT7TiKuydZb7oKPaJGZRz6nC9OodtYttpCj3JrTSR8jP3AXCinXd4Tat6Tws2XxpDXSl/g
7SiwJnLfw6VI4kQuPUUgGnH2rLn9dzMiBpogPGYd3sm913pBiIuk80JjK99IBZqEUR0Cw+4lW8eO
3HfD/JVdAQ9fldx/G2lNBQBKl7ZgkvWV9YslKR5Znru2z3UNKLNqUT4r1dnTdBTS+gwqidORC8ll
peVaKWs+ruw8EqoGlPFxrlWRgZc7LAaLDCcuuEZIulVmo7iTtElrcU20m74hWMKJVLO5eJxJVSd7
WGbMVO4nXRFhabNDSHhjd4p7nsl/mQpXLpqzBPWU+U7sUrEw+kim8J2N0+rpqgQvXfsg3oPLnus7
nrBdAUwnOU9ywczlJxXpXQNJ/10n2hSivdnEn6zhmkmsSqoz/a4qLXw9UUg05P71T2mZMUz4sSg4
Uov/H8VFrB5aLcQ5zNO9+rSLJ1z883LtyuGuALqOFD6JfwBm8kRsCk1X1RxZd42LpwihmoFj9A1q
TwcPfdc27l4+0sTB/YokBAx2lKu/gu9skh9bIwwe4Jq3KrdGA9v/OBIblfY+5uhf3ttrpf7Swc5R
Me3WI7PSpsii5gKM2i4GeN5IW1CKTbFnuAVLmKeiU0wbwtHnrNnbhPBong1PuPQfo0bar2/bRfuV
7Xou4buo7u8ITi+fHQkDVHCyTiL+VKPd+PMQz2d4sAJJtNU5Zl31Ci+IgX45K0lH4vhnSO05VOBv
UmSw/sPvzrDYh/LTUWI99wQLwYOIHwsnls0GahLnZuKsP9niBxSynkxji33AMRzTs0t0hGy7NavW
d0EBDh8+QzCxGKk2+7eqt7G5A8kBdKZXah5DSM2zINZA88kaNllrdw3CYysEQCSjPmD/qKdSG3JO
c6yJmsi0lElocAEO5JTnJ76fXZlv9idXQEstpYRsEtgTCHI2r01rtCyGNdDNjeficD/a38Qbpjdz
w3CJzV3WWNxdordzvHQMF5vKiZz1s9/ogjHsWFiPtK7kCEMRA4m4VGWnxdAkH1TNH0A9HqsPbr7y
La3avchH0zwSUwmbImVEEr8MByYLbLO8MZ31Pc/dJENG+MNV5Rq5uzxlwe06Z9fvwzJBYc8VB9hC
BxLurPIn1gfbKqcwH98wcINL62lfez7MAJY/+UMqhfPmoyOJupGluXsIGh5DIndPifgYRvrbF3Oc
4DzIPOFnjMz6pElhWYaCv76pfNIRhu9iaeq1/YXi12gUwjZU5vFLQJ5EGQV0curPZMCS7g/ZGP7z
5buubn0RvcGsnehEzcjOqalx/zDkZkZnGMWAE+PYDV2xJWAsGrhGhfix8+3QGY3hiGb3Iapituc3
HgSAdVsPEq+ZKK4zQLchmYIEkXuG9vXKwz2L7zqW+yUu9XB2JOELkIQmiMbhWTf2nsCXqxdwFzQQ
svoPxyjbBkG8YKA0kCldNTMoed5RPvcPgn8Iw80Zc5dPeZkrspNM7cVFdB4EuSidWJUfsACg6TEI
svk+5+XsYvWzOXTiI9eZ10eUfCeW9kXZ39VyYDADBV3P2AT068YTPF+mtayAiVxR2X6meXyIWB+u
lgcebwhhGd5XZ9LuCCfZIpgWPInLKsS5KnHORN42lAJbzixrdwoHtZC3FYyVcLPze+h9qH7eXyOB
FCnMMRduHmENkfTmokuwwMS81kTzH948asJB3NOmwBmJHD9xE/L4zYhxqiC5vGamXJOvS+4gJAnH
Wv+9ceWhB5gJwy2eKZOKo8Nvs+Wf465E7L4efQJ9znSfuc0XjfY5CbRZeI8pXmWMVCDCz5jB1e4A
7wjtApdKVWv1mHsUALWJ+kACuW1EFJbMHF0SakfIi4SCUYGr6DdeB5p6ZMSDOSv/jYqNZP9D/4O+
lkGQ40O+xaNHzF2RYWsTCFbd6422S8lK4oIkCqkLRb4H4BQ4ebv0yiZGxLaoofVpiT87HaIqb+4c
b2XSeJiqyXJu6DwHuV6EXB5TgobSoySKiDC+DYRtgoGUfLWCUDihkkXeiQkQzU0dD/tNfJOEQxa/
N3vlitglbxVDrKpMCJvg986Pis7Mkv/lUD0lKGgQ/POhDQa9RwtTc6HINsEURwaZzYXIsaXNCUoo
pe/WsJo98QmtX/qcV+bP1GEM9sFXleHf9HQxCsMsZMqQBKENN+wZV8ghU0r46NgqL37JFZ5aw/3j
2pEYhAfoVCCYvbTxCi94kfQyTEATp2AiwWqBCHYwGxwQQRTe03GlT/JcGOTiT7Yj/EMlQe6c0+YA
1hE4SBSs9dEuGxtF/iIC3x199BsKF4srHZ8q/BrbQ/Ma9KsNUbJCXEP0dVBtA2Khfm/Q512ZFaIa
MFxr70Eo9Fsnrcx3uxiDUwKVNuzxAgF21XXNfsuzIGpGpmYixDJTS6YjR1CFReCgQB8FxRRWDoJy
s2VRu8MT40xYZkzkUd2HHmLiJXqJPo6KYd+cfC3msL5phOYJOT981xGyVUJUo7353EsmCUg7TwwV
V6q9oNpZPhdlz8VVZ+UPVcING1LRt26SlHbFyyTKc6N6PblmKOd2uCOubwSNlI2JE8M93Sh9lPGv
Q265hNwAW5ExAYJi0lGxP1MC6rOZmC3gvJ7cV7WiSB2YRK4A3EH5bir9fdgMv++UsevuWWAEIuQ8
2mAo3RfF1YwA2TKhn8ip3jT+FOwzWy9Q3T0Apz9XATAviYi2iYmz0eyAOrDHMdQYN2htfk9upG1d
H2tGK2YgkPcC4dAf90fUbo8EBWOfY4eugvnPlGPmap7WWD53ZbBc1xPe5pcOscP4GyQ5RDncb0We
DeL6w8xEeCQHkKnJgk4nw+DiWjeijuabp4UkmdUPvPZ8Dyt4vGQqm6Vx7FDoG29C+SKrEZW9G/KJ
Ld0cfD5QY8dKrfQHHTWdWd4StLuuMSbWQCMGyUovPvrNdK4OOh18SRH5RJMU/WYcZOG50x3yLwl6
zPAzDwVJ4WPD6CrYdv7eUWg92JCa6X0XxdXV/mtS6ftqADL0yR4Sql0Khvm6TMGsKI5ZTLyfvgFi
retFoY80I7ZUE3b1WAeuDPFPn89dvsxyD75KSkLeMMLgtSvDJXgE4Oot1PwoWVGxdRxi3SRpxgT3
jKzBnsjSW/wrFiphZVuyqxNUc/jXTTRKvkuX9Wqzt43FWZBUrinZSJgJyn9zk51sUBVoHYZTP6du
Xp+6JX9q764NEseHl6lpDqBeFCxKwpJzrjzErl1kPC2MQ9X8od/BbDNqQ9xMsL0deCdDA2JA++tU
z5b5/8hNk33Npgd2AOXCtHiKeNijFp/Xcu2XroEZqV1KTYxUzqAoGEgrcDm4X/XC8JAMlEkk017H
JdS0TwNgvsIxyT+5mQTiGRd4THbugYbuX6uR6ZT7l6ZwCjfvpYeRnU2dpPAZ7GcvkCYy61LaRO6e
CKcLo/1jh6+y7oYdzmjMSFnVlrzB5w4YreX4IwWAHp3bLBsLeQ4bPaF67BWcLYdS6j7ELqayicZC
WAKnJmFpvA4NjrEie8fQ9BHouTgUix5ceFBYBaY0fzkU5+Hw3PkVr51NcrnHPu9/9gEb4U9s35yL
Z+6F7J2+UM8RaJOgZuTZzmety7agyUXxT1bIxlHXZiSLzghoCk3iWe32AJeBRoQlgQp+qKU7y9Ef
hQYYxv8DmTAD7A2tF0vXPvBKK8zeqlzWWMEqsn/dSz5VN3v6GBSoN0w2e2BnR6uDBWxhag38xbAu
34PBZNd9ZUQGBOhp6P1Ph7bAZjfJuCPdgy2MSXKv8p5AnzpPMXlm3UwY0qJiLirZtrwBny+8p8jd
aEjvLDYy3gsNm1rMeAxUlHVHZ2BpWQTeown877yR3b5XfLG/A7WejWK4HxUa9MKhHyN8kBwx0mpJ
kR2zBYsWS7h65CeXDqujmggP/Hp0o9Avi19YCmD+cePTnPkc1ldZgCAy1qPor9jXEZlZAgtGIRou
CKTQ8Gnw1mM0gWl4a+DYm8BulxBV1BW6Uyv+EeRP9SUJXDaEhqBpGuRfgYq0hGXu20p380W4jsf/
qODBfWbKvSg8ekDijqIKAuQL9Hc6F9FEn5DsrD54C+bNbuYCCJ42DibnWRcjLDLd0myynIVqQsOE
w0srI2m+K+DTinBH/Fs38ci+k0NX4IaI2lVwpV+3sjZnzvR3k6e+4n+gJuZhKYBky5zOsBPfoAfO
KjHuxaxbNkKwENFgQ1/uzvEFgt3mPljzqEbBYzmPaXjQ7Bbp7lF9+WSZyMUG5Xr0D2QWYYhtszbN
8bHbvJDYlnhabkddzUcHBc/+n4DRgI0gYgq7IwlYBYBXeAorZwSBiBsqSTm3rVjsV+pQQGJjXcFU
ZlNhCzi6tCVXyiaXaFfhpeGI6uRdLvtGQHUlzCPDAYh2jqXO9g6l4Rtk2SAaV2ik+yZ8P59w0peG
0WXmIgE0KWGmk15QvzqPEsiYWp6Gc3XnCgZy6AInK4D/9V2J1x6T1t/39FvMjsaIKgQrNE8Oc5ts
qhGKFi3bHIKiIuDL4odB9BgKA3FI+P7vbF1CFDAvSzFnSyOZTRHOqWBc6nPjGj+cfF0EuuZvAhsQ
kJs7kX94jBBknm4G0AgSBmC1ryQauwHbgRajLq4p/TYcVe1GJl6/iHZBtxEYUu+6/+XMIA7eJkky
BqFAyVEJRsZ8StncsyfR3e8nBmyzO339lhUzyjlBJgLlffWPRveU+w71SOUnXUBAbNbAcRmlPBtT
WHyowJioXS8TwwCqO7P1dcIg1QrhgfSqw7mofaY70q2Q70+8Aj1WWuGsuupKGpB0TG0G533CvtGZ
rEsRbXQbOiApeLKypruOChM8qWA9h5YLNgG1FAeTAGKyj75HQ08boo5rImoFLdoq1zIaiTIWJbou
ZVKdVG5LrcJ5L+9gGIl1VXbySZOzlqtjw/ltg2UZfZxmoHEKq07XqRBI4jwOCKnKa6lQYg1EAkDn
zMeZ5+j88BMlTDQRQ6UJnqWKqn7+bmnr8wmUyg4HVfZMvkM5mrWvnEwz4GloBehz8uguKK4SEdg9
C3vVuj+NggLd/zr+f4C0k/rOweuSO3G4igkoukiQE01tnr9EDZu0mAmx62h0FS0mWg9sZAUXs05c
DLbbPBu7Mv5excv7d2YdyhgoRhAocurijpYRZ2r32mnJUNZeGug1IW7U2ps/PK76qXr2BTkosuLS
pJqfvKIyvk221FpZ00lt+76d2EUxBb5oomo3NuhTqO53RckfjM5uvUwFf9DRcBs2kJH2CKEU4bBu
hoyit6iTv0HgG6pUGbgwOr/eTtlZsVIcUrt260qTFububFZX7WolQ/oAOOHaYIR8u7BdeJ5MYRiE
7h5JVB/wBWAftUCzRLsgMv0L32CACu1t/zRcbAjnag6B6M2JSBkq/iUt9DbzgFtbmFTOdmcSkQte
D5095380xESp8n2fQgE43LhjkK59EnQUJv8CvnurECEc2u53O3coGTyZ3FFBj+jau51Lly/ZdUZP
ZJpcvocaH9CDg6g3YDV7Jfbilia29cM7cmD4wIRDB9Pac/eAxZNqOdd8MKHBEaZnQaqH52CzmiFr
AKDLUV31hRDbuMWLQvoowWXL4vxwB0t0nm+tlXlxNp4kAjBvRTpPUo/pOrBTCxNMGJNUAEfObUsL
Y2lCEMzxvZMGr9VitJCpjibhP8vPxwzKwExCMfkK+HYkHoZnIWei2ouCE5OxFaPqhmxB7wDGAxQF
oSNor9olvbef0aRW/Y7rMVjfqUx2RQ+DxMhm1Q0Ded0K1ecAAuCh72OJOT7ftDutfYUdCBDmabQ4
cyTL6i60z4wNZNE0llmXqo2lph5fZq46BFAeDdeLiHluICBcwqq+E6IWkqSeKcv5ESK8Nd+MZNZx
oy5UTVHX7nMiZXpY552npWIE/UPuE6bjnWwoTQo6kuOW+gSulYPl3ca3vky/vP/psix+iIOic1HW
hYiCWMH3gbvZ2rLton3QdYiiGtNKDnnHyFQ75UcViWoPaQZjGQz4GS+swD91rzxVEDX+l5yVhYFT
QgpPBxrJitfTZW8cQrkJDqGCSevJXNz8vnJA2e72UcCz9/VyvVJV7BtmTnNo/cho6IyI1D03174d
mey2xHBVnytUig36A7Qz6m3mX39FgyVNKvf23DQz6KzlsI34lJksZsJBgEip8zDoKhujGLNtn+iI
j3UQY1a2rmPQWCb10xUj5r8OiVOqCmrDJpHM+1CnIf+UyeYKpzcPJfv4n7oyCPbmgSywxK/sFUkP
h8dJEpD70cWyDFbNKpdmxBYfCH2qCn42Sz3QDD3HTXrysZJaWakay7Ln6WVCGlkc5QDxxcjCwr2Y
z72/y98t8mMq67eGbp5TUx7aHKbnNzzTW4DjHzBiyaycarc59c9P0Id0CJAvzCdHFLxwU8HYIl9N
gy5BGsaNp+m1a9zXHsOAVFxpLGz7m+nx/JVQN8CM7dgC3RfFvcx9TPxD5xDo2FhPJCIYP0ddZUkq
0I1HSqUO1TPsPhaJc0PB6IPUyUchLi+O3IC2PihYSS/4/xRRZ8h7lqgNFVcQtrHjzztMWqLvXYd+
Om4mlrlMhzm1AOZQPLO0g6j9q6Fj+GL3VrEHS87XeVfgwwjZZsAifOhK0ofNFQJAxMMgR8ykURxn
FUn6c6x06a/d1Erw48ufITKQ1bAppMlqdrLLbrZqz3Q9hwpmNvFgGNeJOwdTO4iqUfR5FWMX7mIn
lvJ81RaWW/6bzsDomP64DZm+1sS402cASOPIVmLHC8I+1n/+gNFrVa5SJQ9fS8IBbVrMocs7gzSv
iAvCaIX2qR8DGkcD2nD4Wb0v6glwUpySfgv7u1M4xlF+fUfqhXs0VME8Vxe1GuuZ/VVAIJ/+9qpt
DkgkgShpd+2AaC8b47BhDsfSJamY2J+/5yDf8uqYwy6yfN53kC4WqeIQ5zTAKb7TgpXnmiviNwdo
JOxsez/pjbL5DX4Dvi+hCtoMp62e7kR7aza4wleST8bf+PXOaMJ43wxLnKdugYTixQXflboUT721
AGcZCCyDLj28yleTOaAfKzX5vnPoOfHN7ZYuFixXuRabH7OJb026RGKfgNtwpL0eCoLp2Z+LoEt/
1PAHcXjP9ST7UOxOuAl+um/8FCNecUnx6tEQ8wSyn/xlzmpn+lklg7Ya2pXfhh9hs4lOQy+gahW8
7OAszJtjHEMWrchOgPPEbvt5jP5ZLfkYUjXgyuotgPt4GQ4ma55bfuUC3OSX8bD/nDr78wkKxBt9
0JFSkyxWJGBqZxyl8A8BrIx7iuhaj9mfsF2JexeOMW+EU2s2vhkGWJiWK4J1eSmzKtQnI3jeJKjM
8dvvxapeIwjMSs338IJdVdMQQ7STq6vl84moMwLGBDKx4niVRsNHrZRq23nSwMaiCmsWpNAevxya
7a4cg2zoRLwdhktW8j1UhQlKqzoTLLKb0BTBYDfG+BVfPo5iXTedqJm1UdsRIfFVNKaFREat+yEe
ttj7OLI+r6l96sdImi6Wf57xd8rnkT3e9mWeV+8Qpj+hIeZX1I+BdY10G8YWuRBITADujfVetmmJ
gVa2Vt5ARA6OkZySurEe4Q57VBxjsXVD2yXE/JN3kJLjEw+EM1or4F115pG8Ifa6hYdvZQ0VXxdB
zzk2C8a7H6HJYYOqO0i681ZjUQop+2K2TLXSAmY7kCmpuI5/vz1cjrY1iRL5XkS5POHkR4yVK/F1
thkCuzvt4hQi36V6ePjEPKARY6R1q9Y3e4xMByZSaUJ+vM6UwtTOpE1m/daQlHGbu3WUCZLu4/Jv
WfVLBQGdAhNHNXbGCicc/Amomm0rYJfaRHVvyKZsZBuGY1hO3mXRedU0ZgqJwjgzBKDybaAUML4y
RMfIo10PU5Hn7SJ4FM+zdtmL3b/o2+C12yj+VyMseb8sgLRyvCnm2PUh1Muz814lO1qv8kO6vfpV
9jDxBtyRJAxc6YAaOvKwG14eBgWCZJ0U1ZgOT6MfgpJ9BMkTBfPlLi83tRt+gX+4jxpu1Z9l5n0+
F1fz9LJeaHDo+4l6A7qRj5Z5l/JomatJ1bGZ6plFJ9zvC8MqVWg32bWl+R5p1UsKRnhb2HhWTXhO
4k8Nq2W0NdpsR3lrjWJZS62q4X8cxnygfj7ul9aDyvQZM4vCxVnbfIdhovzkEufxUyIHxUGrjewu
lmIyyieNw3EdQPUhfqzC3olQH3eg19Hhzz0BtJvfEg38+9ualThiay2/Pjp4PniEPRgNADv9xPQA
SZW3biekG+Qt/qm7nZpHEqhmFenh5JqS3/wtT/hO987YwtA7E9MZzfQS9Wal3rkBnL8WfTzKuAjG
Y2/ZdSYuNGOC+9q6/fRaWDSR5kRSlk0MQlVQMmHSjxUyYowu3TcCN0qZyPsHdKriFFbsQ1NkuAtt
6ecbtCgypXMM/01EPL923f4bZrPUbgRnI42RfysedLQgsk7KFpwH5mZiQHcx6fDSpsq+eO6j6EmH
1GoO/0ncfkRPqDszdoGlpy8qCyvnj0trXjUsAv+iKg4XUW9ndyMrG83VWjRmr+VTTkduns1G6Yeh
/NYRxYnZjiANA0HSOtHfu3ncLrF9htiM5OOtIIwt2tBv13D2Bft56c40xEIFLhNIshT3PvipeSGj
S37h6xDbeVPCBEscXFZWG6C+48cNvmr+S1WRdYnVz8uld4XX77V5Zkt+8atbiaBW+YXi9OiCZCUN
KWipcR3nr4FWSopm0nYU+4dJK5X2tTTHnc5MTtRW3vbC7EtJ0MNAJq37kvy/r2KsQCPfqdE/Zev6
j9/aZMQnN3G2AHe3FIcWoFQjQ+3lou8UlIAKn4m/HRZyFIaHUdGrorEYZrdFRvkGPHplpA2gR95k
nEfU8IeL/wPrqbDXKWPMFEEKGAxOWrvNWtF7ZTdNLCcZnKBwGWBCUYNztzPdsoCLqKXnEnle36Fx
7jXWosJ9gMzhJ9fDs9f3AhlVTiicQYuNPjwb5oGw173k2uo4eQEZIBu1gADsZMtYOzRavKQtoaIh
3bNfrAQYOIDktHITGRmHk7CPF+/vh90ovcAIt8vL1w0lMmQpk3ow7CLrke/xKjM9mthvRrJxAP2m
prdnhZj6zO13hzowa6cDNmglmSE6FuzEDcKkq6ASrDvqloZVYffyjZljvlgziWEjREIUPw5HJQZG
6uc5jzItw6TWuPGMP+gWdIjmm+qYlH9lQ+O/nhichEx/2XinNxSHPi3IsT0uiJ4MsMk4zSI1JnCl
zjLzI/jOIvhJt3cMoyUd18N7UDQ4WZ2FVRtECeXmHKhbcE9psI/nS9f9RGdWd9XSJLz72R/uVfgg
BSpZQVkal2Ld2wNCpdZT1/nzGlBFsjjsvpjg3vKEL50ksLSb07xk6MeJzxyEe/f6y3xXnJq2/4tO
9XYc/phIx0Y8TEAsjttFW+Bw36TIz2fej/dm1vseAM2nJX166NiWKqw9C9Glb7ss+J/Wwh+Ynujl
01V33ZMTYdC8qcpT4kFP7zggstLyxoWHP9qn6jHvD3KtYed+kl5yhFGhRpRmjh5oZYp/eRJBN5Al
pJ4JB6Bw2Ta2klq+w7Bt8Rj47mT69NiLg7rLUYj1a6oIoo3JZsswOcaL94lHRHjDVA6hOQ6cggUQ
FEwY25kSxje5aIR7N4Vki11IPs/b+gCHWouPys814Cx7xjm7jKmYcrZMw8PI/9HvCPY5dH5yQzSG
N7JnEqqZpFts8VhF2E/zTTVwA+NENSkVlfdmFAtuV2vtnLzKdp8koKPYN84Jf2iMszARLHHApETE
7VVl1U35dXJClSz/b5jTA46X04urdEBSYXqIBN6mWbEunD0jvraWDBfrw2Xu6rCzlbJMwThhIzNL
Zl99wa+dTclyxdEsFvrMHARQ7WKaJdbSBikx3KEMrperb3wwJUxjTZ0NrfYHEiAFKLd4FJugJIPb
Tb6htV9tfahFvVna/CkZHAmbybD4ZhJbKKsFZBX/I0hB2X0JYp0TcwOl3u9CpiGrPTmH5mQB+g7B
gloUn1yQoliozllnLpxiKKSLa0nQz0QSF96GRdlChuPScMuz6DQRUs8Ax9BBrg2cHlx3+UeVXvPl
7xZzS9y5cP2xgu9o04IyM3NJyDu4peMHfL8AM2i37Pqhhy/Ql/CSoCarSIy+yMoTBbOUxZEdFDCp
SBKO7x9Kj9pBwk1D1ecT/T9aaCZD5X0WFSbTFswhegq73xWn3gyWEf+rHuIZeseiJjyY5r2vDQLf
Or8NlyK/ULNDjDlMb6jZi04Rlc/61MGb/CrBBtvVFx20hpOnWW6Z9W2C/NMMtTos0m8tK8fTQB6q
nr5ll4L1U1WBhOGqOOmsn0mr0tYmHqVfotKoOAY7HQxXYYaNKjGKDrWbH+tPlP22KIYNoA3mCepi
7Jcfu8jCRUYbF6ue8InWM+GRVBqCNQ5mtXV70KJvuIC9HCnYgiheMquLCpA8HfjKSCzaAC6kM6gH
Lm0Uws7L2SakGPSU7F7JGDWQN/QcMEu9Dc25+WqUpFDCyXEUWBBKJk+Co0HbOuuFgub5yNNnbBu+
ObufQQl6QxybAo49Txn9q0wyxYVwNU2yxej5xcB7LEXJqHYSVxCTyogazG3mXGAt6D8uDIiNzHbh
6SF9yK5vz7hZQlfXWKsYo4PbUji9vZkDzQvy64i5prN0FN2cXdVZiMaTcIRdYu5tqcFkwLJqgJHO
cc3o7d87wUoN/JpQy49T8vikQGNVgHYK726eSRgIUADigkUEmtoXv4I0cbplMhrmQGLWnS64xyyT
uAQA9HJx51eJhb5A8XJfyRT5/acHVKRooibNNUPhDMNDS5+14AIDQuvvcW3rHWly81o6TD9MHGJM
ESciopxWDEym4+F4O3zPziD+9BJ0TOBYEZ+9gAAH/qkE7m5fcIuKC5uG+9+GAJG9Tb3/e3WKGaC2
3c5JXsx9bYUlUaTu4a4g74Tw7+wxznz1bUgJD5bFW+EM9Ior6w6FHFZ6oC4LOnUfO7XwsdnoQTTP
s0O09I/iviqn07RmaveRUaCDMD91jL4MQgTG0WlUWcbddtuxaEkK/V6Np/zDquS7tS67ZF4HOYrT
oGZubWZ/vvHYP/iHou2Sw2O0zc91OTLtsuxQLh45W/jn6/NjXrFv7RKUWFGMYRKWic/25THo6UF4
1LYvJYY7+TC871fnUiB2uE6qvspVVVKNqPCsKVb3Ic3CSJl5vHt9Z4RoFDkcdtzsc1pLRiIM1Mze
Dm21AVxs5BTj8dD3ePcbt2MXYIziFqYLDqhElssD6Bd0lcui9Nsw61nB/sVn0uK/vi4k6PTmKF7O
6J9JHnBgiolEROYlsgOuFEW7PqbKuoON1vMDbir9GM0zjIsYuB6FIuZYtWOV9bjVUhNplHwk5lkI
+fxGiTM16qafOInF8BE5/6K12UQmBC10EhnUBYa82rj4Q7Q9oiUbjVqa8R9zM9lCVTk67DyqqgZo
YWWtYWVgQqjiHRVuPZJT00lxBZxqOLv7JgO/Vj9lTgfPAsgrHrYnF2EZfS6AZVDLDEasu/iVfto3
ZUO3klb67/rAmbwisMGMKG/stdF8vfkxw3YEj5acn3j+PkDmyFcoWyIaLH44iG4++/58W9hzjwfi
k+H2VsHoxoBDMsPLyg3G/6qY7599nCrRa2827JXGxtYz1ZX2XgQn1nde7Ckh/kZvmAGNkCNlsyGU
Y+V0tQ/yhV+I6Nixn7PQgRhis7SsSiZELiI5jD7b7hx+5PL5hl3zFJGQGicO6CR8nNWtOF/Udpvn
9m25pi/mR0r4ZNJw0yx5Ll2Ei8gn/Q0TaTehWowxinOjoA95okjRmoh1uQuKMfkLlGaQWTXm6clb
QxIxDCn//JmHvexJXfilyS3vR/17ZGsf5CguLPNMqAFQhrkyCKeb0PkCaaG90Tv2GSQX0mT9TjaI
zmNfWs9V3BSupJAYdcxn+3Fw1TgwMjPqcZtNQRVSXJ5Se/erQ2naHaJmxgyuc4Wq+dURD0BsCKzM
fbrcxLm6+o2Z4llAkwOWO6Itzgz40U7JujWcUiM32uT9fIvSW/NjXL1GfORUDylK+W+yvfFv42jf
XRgNlihKu69LAXpavQn/op6dP/q9o9RwL4dEeHtC3HoNzVzTX3+In+AKVwmqNvOShfn4pv47ok/C
rz/MmQLTbIo0OBms0JmyyNvjnJtopLfmxKagCCbuG5nnj7H+qWNAEV2YdNfPAzButx28RzRrCk6Q
q/BqOXBwivqftIhK4ZQ2MC+MMGsBRVh8Y7h2F9NX+LVbDm+qzTtry1ZdeOcKXThUd8E3hBpvBWKV
9AwS+gzRFltb7Bso1dZoFkS+sxt0A1j7SzPUi3KNpW+ARPvieIcboZ1EGlSTuvMqn77lTCmMFSIW
cKqGfPCzYs0XdAG+LbGVSitjS0Ahz9yVIS84gwjj60lm5GAfi3csMwuFzGD6vZsYL3kdVXlNCOP2
rtTolcMGfmKB6OFpqXivz8O5wQ9wjRXZmDsZHy23yUCeB73kawP+t2B1sezqnfBQiZCWSWjotKn4
IURgC8XguP99bIbj+N/rUWb2QLQpt1EVqyJH2CIx/LZyKe5xdctg8N0m05THsEc8Xswqep/YVxia
e4i4RoscwF5F11JEQpzOmRlftotbVtvcbJTGHx2UTRukkSQU/wnkRBw50EfkDxP4yIoKOlRYTjD4
id+M9VSCVkKH0wrC2+ahuf9VSWMCx6nmgu9kuRU/ZsXSGd0Tp2BJlEF5crDlW17dUJTCUDMm4uUy
ckipxEzVB+6KpCddZLgy69zvMA2CEPncqvZF+LcvmViYmiUJ0xI8Ve3uh3MRnfvHFDE45brxPYnw
9BLTptsoN+uT+S06kbbwcsBTPe6TGhOkbasI9Cj3LyItjyHPLt5xUz4AdpL5xOmcq/VFDqBiM+KO
SgZCPTlRhRipLtz5fDD2bKXEPzKNnc4/9N2pRILNeQi3pN4XNNmkf7oHwUNchV/vFAdtBO+VCy4l
b6Tjf/wybZA2ZGw/wGxatkUUdnOENSSdIC8PN7cfX2TII+ZLXGXsApuEeZ9IaiXHwXyPehwOEh7p
HELfRKZdsdz0jrKbGWYTB5XqjKRC/fCiH5H7T6Jbccby3WlLfvMSHdjikk6uRZs9zEyFq8ALIY1S
18UAAzE/DHJeecL3rMpAaXlAXf8mwksHcQ0f4HxOzxRmEV3hJT4qT14aCkAwwJWv7+W5XbqUG9YC
MWNYUIUHsZxHtMThemt9o74gNor7NvU3tPC05Ol9kHZITidHtnGm5Pg/dUqSd8VIpHnRHjx3ZXcT
dPJr7B6c0zKNaWjgDJ0N82/mj3W8FdmGe3Uzy5rjA45I8vew4a2ZqhUKTfGy50xQAalXWNZK4KQ+
uduMNgintuKPwSUOQdSX4hAWw/+HtoDVckqtqUf5eZC8g84zFeqlONuLGIMeD5MuEp5QXP9xr7Tx
YFX5xa2khkErOak/EOl867Xv4D9qW6lWN/kxdAHGq9r4xqsnnvETkrnOOu7OAbcZZorxK/VlPm0W
bcaMa9S0QWdJdgs1JhGqvi59pF3/2jXGsPOowIXR1XX87B8GoHi7rfp0urQV77U36sjfomZzn2AM
8XLWLx71pQQ51oST9HlofC0zEBJv4KVpwSKgh1qxK34am990aJYtcFOLDACUYmD4R5+brhVZ0BQs
/epnIp948oqTIAmGLvZGP3Qk5uiYJr7BT9FG02M/hUpYRJl9yVLE1wfjiVUeCQSqk2no0YmfaFLz
IEgWzXxqYmJYfgzGDVwhkPCtqAYauxLRXpeUqsN5J6EUI85pdHnCHg/DTLwu7z9Qyfk0HBPOuDAZ
tdW38iSiSQjApvuawfrz4s7swZlY6m/ZEIcJOQUshuqIqrol6Xf/ILM3psByjelbOocJGYuSDcyS
oUfSy+hlvmSjxvazFQAJzKxZ39l7KHHc7AlzQ64Wk6Ms/fPbAGGHyind0BLWjTy8khP8rup5fzHz
9pvDF4JeDhWPkOGu9KKhkTT1OU/x1fstxuJbps4If6NlYEm/32mI/HtZtd4UCcc8O1PCte4d5nQo
7cZ5JN4XJFfImaIyVSivtcrIzZ9IVmLUYgeIxRG1kjqAni7K+oXnwtvxwQ0NMI6vC76wQpKK54zT
1/Q9ttNxfcYC7hXXASW55XTKZjKv2pUbBcKVm/p/3XLimYxofKZf8Xjd8e2tEHYx6n6S92pV147F
h6xRx2JK4RlkobUS7ICJ9RN4ViuWWjKQQpHCLl0hnP4+9K9vBjS7OZJ5AuXY01D/fvECTKYNCa2U
C5f5/l3lHBwQAVLRrM4H8BCH5GWHf0bReSzL1PRSe7NiS6QrxKXl51y/BzYQP8oNV9yXXO4c5IUR
W9y4dUOpG5pf4SAZDp5UPkrj0MIaek802gmuF6jgxjH2mqaEN01vHarLjPy+7GsNUI1XUf8/X3QU
QHPEkRWG/JtKMNBdZ4pkwyaD4HCDUKhlUDRiDBYzt9CM51Xidm61de9RHQ4O7Oz4+5/FzHo/0i5M
9btQkhf2xupybhOg29cal4Ur/e9poSbdy123J6+JEe0NevP5ZQbCMd/9krBRSGwZb5nHWFe9Yavr
COhfiEP2D/LzLw+4fO8Z2lNG8x8yT4SkbMlCpYUwpHd2L95DVeyLZb3OtGRIE2dbkbmGegre9YwC
KoqK2KJKQqxtIi+MPPAN90NoiAWraorhBBjQ9OFwLgP/Rk2xqIMk6XOX9KDft5p8EypHKBOeSSDn
PcsyQD0/OGgzQOnFH6PhTt1Cgb88GhYF3UakMEQ/WtijWXDTIu/1MRWMZnGlogqZg5ABZxfHT2Ug
Y4aOS7YqRJ55Npg3hjCcCRYp9g2lc6+MorLgGgca7tuGx2l9WgF4pFwWYzgi/5UeBH0sSTjHvaEK
DG2pJh1MHYOYRMDUmVywsjUezQxeX82PnUksWx9CFNEL1/zbProqDyjsRC6XO+Dgpd2r7ov4MhPK
ykPocgAC0VUGCJhqsNg5JktKh7u6b16Rv3Hl7LP5OPrwawl0YQNO+iDM9wZ3aXrHdbTBB024phB4
RR54NVpExv4FVErhR+INcttJp+CWO5SF9z/GDH5aeTSZ4Ws+USFPxcvoaGu9JQ/KzOK+g7fRa3Oj
pnmX9lGAPp8gWTion1bEoxN+e0Y2N+64SC2uhLP4hR8kuyiVp6Zy2H/3gFz7HfBKsZq8noLZOG8y
Z4WdbXkY1hqJ0zsF8chSvQ91pR0yQgMc6UpwO9yMdywVI7ePQkfG0agFUZinDV5mXkSpS0nUlH9u
MqwTEsFY5hWlGEtOLfJfvmcrKQ6nRMyb2eJlo2uDVt0e6ICJ9zP60luio3Zu8cDkRIggxuuPdtMl
7b5d1UkEOCjyQsB+RnZfDNv3ftvfIKJXYZpkhDWydF0+SVxrPAH2a40In2pD4/YeMB7FIUyvCEHe
l1hZkkYO0Xc8av4U+5vsGbvKCGkHQrWwONYw/ZDG+NL58s2ZVYrAcwmQjaf/9fdD5SuRlXo97ozW
3kJLwvTr8kS1TwJLh6GRy+AlIpkFZcpB/LuyI4HWFszN5A6vqBnE+x9iHepahtYN2ynzxg99Lc32
DsJaAhfP+rBQUapGAz06bX8XoIx8W8x/1FOkv0jpemCUOF/LHzCqTbVfcszdLzubOF86H294NXrG
RvTZThT0V4DvnFK5T4MoervSkEQilmS9x1YGTXjGkZfVgj2y7DQEUh1dK9J9qfDDdAxX/iB7fpM2
JI6RUIwaNCD5EGLmixjWvFVHNT3gQLdMFUv0CQEsz/UGO3Nb1ZRgachgRpns9agS9HFmS2UIV7tC
G2lkP+aJPzAI17EfmX5oM+GLLvf6YHjpf7JL+VMs6wMxqB+91wWrn5wLn1uyzTOZuDF9iFG0WCMm
gYle2mzmucEYHI9wLNTibbuHBidnNTGqu/3YuV9DvSN3kl8hSuYNbbnmy0anxMyCEV2MuPVqAfrN
8ZjGYWnXEUyf7MQe4LBTsnB67tQLILU+cnXZ93gQG4ZwcGhkXB3uYJg5sxTottOpCp8mSqOv/GtL
miXg9locHj4oebwi0cKbkI+r0CAe00E4Abc+bN5GZ6b7/B8Le9q5AnvTH2rGBQm944A26r9RTFVe
dfoGzTWrsJcjxW4J6mbB00XRwX0o37T1zayqdX69gRVfplJjel+1jjtuyC5Nzl9K3j7qrQne2dC4
qRjWOPmjGtSZOpKY5LRM33rgmsDDzjOVW1eN4cYo7R2+b0ty/Lkw/hvgrxXeipcRqzbKBetScqr9
Hq85ykTRnMw4Eqw/qebuXSqA9+fODPTL/zEKBZDSha7lH9JwD63GTMLW+17amJBcl6yEldE/K1lv
CnsLHVMTFzt4PlKaBGXMjcvEWDXpOmr1iclboPVBshkRbsSCZLEniEeyKqzP1d5CfzB7HoOB3q0Q
whY/D4HqIxPGUELiFavBKP2qD8/c4GFaFx+pAfIeagoMFdTF2Jdd8OFD/j9piS/eTk0iCATQRgDH
pkkycsT6N62R0xFVgNUIbjd4bnShmKN6C764l2xgSNLGG3Qbyd2cIPHGh8YzWmReAZCnoRZeLjbs
Qv9D/jmLiCas8zgLzNcxYoOrDUbISolK5YKHy2VKWAiTCee9tzovDL+HYOxWKFNUwjfrnyb97c7u
/ReXCes9Eu90FZA5cfUcH+82TRiYL6yUBUSUiz65RQGv24NOFm+7QhphnEWIY4Ox9gNmhVbqfKG+
1Qv+uM+S1+pC93IVLg5T+S4tg0Vu1VuqDH8s2SffjIWUD8/g9E1XZqwMji9TQUqPjBZa406HnNQ5
pLBxQ3ERLN3NH8cCSFpLe3R4r6xqwMLBt26ywq0ZpTDeXyZSo9NMCQmvnelPh/y9n4KlHYgxewAs
dnl2kplneNQ6Lymghw5C6fP4B2FVowHJwYV4LtHu4oExycpDMuKAAQak+leI8exfDwkSvdQ88xGR
lLUE7zRB3M6AD1R42y12rbRl8f/Gl0c9f+4PFYDYcU6jaj3dG0BuTOEBDhv/PD4xrB1oVo19Vgd1
rV/kW4wCvY3uMWsBScQljvcdZR9W0peLVSSu66XX/V/tSMtJVLb8wiisDTsTXkTg2az8n5alDgQV
M0teAZAwZpZ2MDbjb0qGHUeceeooN3Xrf9CXSKYj/eev4VLAgMRErO8+j1nv9EmPbWoGVomUisDL
Bzsp5bekKP6hgmKgpGFfalx4anIoJArJXZhjM5zaYNpWKbfnlwwhr0gCZ566zh5rVRwPYflh9KFE
RsjNRC0pdid8tLF3vO5jouaH+9kWvARzDBFgYZKijttkiyADMY0MyogrMGVwkBIw4q8bmpGwoAkv
ED4Lk6boeA9MoXUlKWJIgp5j6IbGViJIhCj+nufAGyG0rn4ZuLHugGXTQI7LDtheVYSgY5g2FNz/
f8ufKzQHSBEKF8xIDKcjZin6/iVomvQcBRtm17Ma4wjNhxKQ32wHn1XDC988v574yMwoVzvtM3yy
SYr4SWFtnSeolpEirQFZBvaGRYO9iVwlZbCzAJbR+L2Cu4USSK0jn+IIvafdIIk4pgMDo4jmXRdl
ZVDgou2Zvd3nsHxijHSJmuH6BeDgC0Tki66Mbt248Dm0DNFrpylR6KaWsLOFrGQunuOR7E5Bs3sh
KccU6vLHBuw1q/fKeGPX9cRfBAtFW1l1nd93HzTleY6RfCoLhmVdtQ4yifpoQOptc4Kk4BvGzlU+
pc5NVibhSMqXWDLC7G3hfBJ0VF8KCAC/30Wsmhv5aXSQiyEj5+YUj7435rBKUCSMx8fr2lKO3xW2
J5N7yMqO3FProSS8rkCMdduzK10qaPRI4+0xpfGwmogeKQlEDiNbiemlf6SwB/MA3BPdbcvsMAX7
TbkKSHukYmhONlQjQ6kzk0rGVV9p4auGnlgBIliFxtnLp8+i+F7C2n2BNwz856e3R22u0pb0j/RY
+Ze/vmppLBgVdUWkYS6jgt2BJMVHV8lAVRMI5HstvB/vYvaFYb04roHzW9sK6C/9qjQlJuwLnk9t
FRuJNL7fLS8NRJ1j0/bFBCavkyh1tqWo44z8CXGEO7w5YSDEoePxBc55tMgEAoXS7varL3Yris1n
tRY8dMNTOszxwuHKJrgyRGs3qKLtMtVZelQgQiwQgWHdB8fBeqs+YVYw/d25N4ca5pdu06r8ko+7
EaZD0el5uPQfMGpw6w6SaVKIZbQAxaSX+eT4zVj0FkrdxJfWsnNx9DX2YY/ekPIJa3D1aoG+2/iO
EgWpJHiDrA6mlJzMtVKqxGurIN0DvUZD6JzUHnYNZZkZ4blmynA6RRgLX7ZGbgOvkPwPHUHeMWgt
14cHeBZ+ZFCVwmuRjIIXMuM5sVmgBLdHql3BjbB1LbZP3IeI31uTEWHD2TQuqHWomacHJJpGb26c
YbYzCdxAPh8WRyc7miRBk0YG9vRiiTs7lf0JzU709H4FUgmTLeg7j3NRP3w9FZf2GZqClR+yzUmP
ysnWH0LAUNWf1IVPwEkp83fa93vuh3fLE1D/0ZNJR5AmrbdBC5sYwR7bBa2GHYAKWmKJ3EiWakb/
UCD5AHtJ8yAJWQS3Qr6ngSSZpL6MF+uYAvA6VOwT2f1VhKi/GIaFwmIh4KJBpZrK7kpikFXHDDp0
FbwbbHX9MtVCH4VVfzQj+fm41vh4/mN3O/QslAoQxmcfyf5MJCk8XjX8eUvVM2A3WqgrV51XOpXf
yFQacprYtpfUxKUQ5EdBmiSPH8zEbbsBd9HPxdn/nS2uZ8LV4bHoUFTJBZKsKXT5nEhaxx0iY7jJ
3kT3fVgrkS4JfRYFbacKZ3jKRqqNBSj2jGyLIrGssy4kE3iuaWEyU0u5Akrs0/LDghDp9wrP+tyt
S/3vq/Gb5INWNOHeM74mHU7Q+16d+DitGns6iu+c2bttz/37KS6phOl2V5sjiPGQgE7766SNCEn2
RvnVJIJoy087ctutkf1auZvcy/846tNQxCOWwO0qPTAVTuAaOgxrqLANB3tzTuSykYvFfH3nM+W3
Pw7kjxKFyWH2AhrFjUgsVGa/Zu3Vf3bF392+MN+4BsCCzlzjDqQARvIQeFh43kba4UjtS5jznLSN
qhNgcLLid975X6Nt1fT06HiXWUWiVUidJof+rIbmK4awURhSens5knf6Em2tMLprlogtk++wOF9I
qwo0LrMlNC+1rEwnKM6WECsHH40DjnOXmt6M3PwyVIbpgAlJGechRgKQMGfZmMS0ZuO1uRTjbmOz
xd8ySXesHN2NzXuxay4Rjl0c9lgFZPPT3BEhzF1zke0NsQ/d1VFTVVYn+1Lmbde/MiEZ0a3edO2w
70deSdOrkIIYP5dY4qo2E0dKELYkVcs69XnfrWdYlmNQev9g8WP5yikknwLMKt2qHK+F9754fm11
p/P+7ppncgeGwts8Crh5SsK8W4Vvq/rGqgD6AL3kFV0cOtIiH6myuAD66RJeJwSrSI+34jjSW+Or
wxAXukUxDJ9t9qLSWoE8TcREnkDEwZ9sRnvDO1PJRCxQMHTdNKHX/SaGn2LSndgAdJhNOIbT6SNH
ADK7/3EKSTbpuAk1vHcuIMDFoO6iuPBBZLE9xQLZeeujLOHC3K+ksg7cGm96RY7yyvkH0dueix9t
6FYcHNJOQ7YvY/U4C7rhNn/yxb6LiC2a98sr10q+2JXwfY0BNBZ8Bwv649xj2LH+3OtZuuwPdnQB
4GA4HYWAcCB3gf7KOzb6u/7nE0sa5PDeIWYtkx2QndnxZI4oISCmmdbMXQr3e8cUz1QVxT0C1Zn4
5HSBcdD5IyaC/dFL5zsakwaS4YULJ6SUURAqYVd53ygDHx1HGo+zdeTFt3QUSmDGNGlkmQUQ1F67
3pMZWXSr9zATx3EUy6lTgZ8Zr0tXSejr7faBo2VxjbozEGZ86ZLxFJqT+6sKU2BOaxZIdIMmFUZd
6H8HeVAC+GqnOqmT8DilJNbvqX61Pgb2yinpQY8KqyV4VBRIpiYWWM/QEeo9a0yPn1th8BQE/w6u
bL2Ay5p3eqjT50YLThpHirVebPQavqumQOzKVov6/ylSKiSfGwQWIyWM2aIaBi5nJ4Lnw2M05vr1
luGK56Hvv76JSJ6eTdHeID5a/XX55auqI25k2P3PX4Whie7Dsl9IL2ZCCuj+Qd2ALNmMor0/IA0d
lAJ9EFIyuZiOGl4D+cBsjFyugGEKATOfXlhi/H0BalbbMFmUchZ/7oeRRczV1TCv1WwHXx6fkMn1
6r/6QMLYJMRnmxsRvszwtvGUTHdRSVeJvajr1u0jSBvk/D5z/QcEbrfJrLx9LqhLWqkbRfrmFWu2
yU2HrDBxfLZBFrPLTWJDKIdOYv73oCX7obgm15mqN9JxepeBbTvEXlCSwkhyfiHDvFM4F8ETIZoi
1elKS2oQ78dPD3kRLHzT9JBUUs94iHh7+MBtGPE0z1NlIZ9IFTpdxRMwKqj4k4cITOkL+0xQuIMa
IdjDkYjntU6k2E7sgOIV2P1m5EJoFWOyawAYUcGt9JyMgyORa5J+WevRzY4HGCnil8OcS1Tx2iX9
WBvK5MbftagRXohMMA4yabQT7c72LSI0YzXO0mVP+ROd9hTrxCyrXBeGCwf+hfcQwa0/yRhehp8y
1OXmMkqwKUnst6bXXxYA5GwAeTAO++UVaZcZcp5lT82chCKljHyFSvdlrtAtnBsXgSfn8FIcEKc8
j9ioOXCrWauZzPPcFQcXp9B3AnQqypiN2BxOLtc6YjVV5FNFg8h0royYjZ/ksE6SGmAMdnDv3/9i
q1cD7pXBVa3K3LqlFo8UY4OxT6u5OHuFCRMDgJioN35ZNMKs0uU72Su3KEGhBgUEu8FkSE4EYb8c
PFc01WxHVb15kJ+yxxGpGy+a7VbDyXP7LdneTiCKx69VW9R8yUu/XHakBOzSuk9PbrNQ8i0JhHxT
fRKZHdQmMKuizokk++Y/GbBqrlPwCH4UGFhn7NSXEl1yvY3l3ldvjVgTTYS2x7Bk9rRTpRLzpfAE
GBecg/+fC9WOTNme6rCDB8LsJ6g21bnyInS773dzODh+dswC9VwFGuOTCoReg3dV4a/+/u3ebSce
mJ6/LoJdk+/NCUFO+B6775E6JMlOP9MxHs4T9mvaUrpbjHoTbPhpYLGWFmKWkrE01/qa9RB/419a
ZjaCiUA2ILel7GITdxUmJZ9mRArRqO01yn3r6J/l8o+TNpfLPQk/CFgGOQYwAOVq+otYwCBOTQ+S
ME8W5c9MUBWUvUxfikilxcZT1SICkPPQR1PWqysS+kJPdc4Jr+swxCiNXJ0KklzI/d4GEGmpmsyn
dfJw9gXUW96FWvvBGjgaFvAmOjgEEbP/OGcI060Qr0ASLX5HH1VbqRSNQBjBhiAVUtkBj9WUFCSE
n11d3QzOTu6YwxtqC8Q0hq8E1svWmfZbkb7YxOAFPyQntfffSQrO6wEyUea/zmqrUDRnbJRW3n96
aiWAlB7t0sYJWsTL79+5GPMbjMWHHBLRGxRuWzlswFVFCJM2KADGoLnvR3caAddGZUrgByP5Gys5
S/7eHiUfTng6cCjRq0R/+qkdOP/9rerJffcNnNFzAEoJzgw78NpiVA+QSUC+hHDYj/4LVQw4PIW1
A4ancvqBQYT0L2cgV6tya2cmb6W5zmAncx753jhUWoub0eQHPWEhlzgmN/MnkXthRv6EB/VZNrOh
DCdTCn4oLlq11YvEGUffQyi7Ca6o+qVklfWZsGOePzUUqM2YL380bZQRbLotcHRevPUuNutJDYDT
Bq8B7COvnZqExrvWJlKJH6VoN5cnE03tcCEAxUloO/1052hbAckMjwAvPD4qaiIFdEtXSQoSSfJQ
FlcRXQ4Dxjrg/+kjr/2NXmqYfcB1aEKCma+SmL6SxYttpJapBQJCvktOGB6xfsqhxEteGqyBiReE
YaOR1ZWUuDmcF/OWZP3qajeaMhY1J602unWE80oLivlsFo1PY4DUnxnV62WjN/b0LI6yF11sGeBh
KE7MyCgPG/GBN3byF/G5S9had+uvreUqidnOq8tAj0ce0E2WX09kKQShoh9IkUy0QJpbV0fOzVU2
8CJBXZbL0myTZ2n6wTcBBjIwqAK7TDsG0r8ZZY4/BX5FyDf9xSxsm6ZaKdEl+hnDZWJCfwj5AZ6g
ejLN6gu4sGxysm5/3bLHOMJhWAzcxYEt3NPVKH3MslHXhE7wkf41joArw/BfdSIbvzU1NPm3eIpT
tqoSEQcRpmTYWLxmJitTAxYxuUh1EgW98DDx3G400+qrKrN4ujDXEyGOedSwJhkwJDohFwVEDkg7
A38ZTrat+6uC0ygi8Mc5WbghHOlYMZN0EZMO661isxpiwGdG33Ows3gFbyiwn15eSpBX+ogGd652
f2Iamj083APi6Bjg9cVAoExP+iMuRZaTuWsMYLURfQenJUbTk7V5LM6pVSNHf9W4u62kn+1Lgohh
3ZlhLiRFilcgyFt7g/u0mTBsxcOy31R4cmsMNOlkiCD9FAH4kLeQM5ZAB1T0Ak0c07w7EPIBpLop
lxBoJoGafg3mNVN+FTTbz6kjnKpQMYxHQ8uADfG2yiyAsV6CRyYMSwyIJdocZgzD3+NBA7Yx0SXL
scalaFGf9j//c0Xp3k5X7sqpCDAzO+pUwiDpsnw1Scopf/MM/3tyP25S4J2iYcZpHLQmcj1Lj/Fz
X8ngYVy6EXMWBgY1Noomq90fIdX+UL00lihJvjGKg14fXcM4T17uC07QuFtQ2t0DbvGxl53fPFst
fW9x099ajgYYsgtZOWW6+8QRkww33Z9Uryv8f5+CSNrmA82gsUhaXL0CpZ+1xoCuSTP4JrntZj4I
vmz3Vd2/tlzt1Yv0GVbHlEgH9CicM+OHuZaLAArKf6KCXbC9/nXu6lsmG7k6XaoVRS3xv501Rh/R
DUImjApihGhzxygjTgD7l0CuKvhvMQCowjQ84xQIrJQVaAk/Y4sX11VO4JRBL/DeypeSOtRlJEqR
saP7ZBWu5L0kY5mdbCi6Hfp0sz1hbuimUexcEocdPqWiz9lUnrj1saaDEl6oLh8phqtgAkAb57H6
bB8aA0x/b71evUQaOXrxeKU4C0Lfo/kYevcMk1+HB7v3X2nuENYIcSGfeTJhj5bRZzAMYWn3l8jZ
NeRa8tdvdxMlIJYAp94qtFnXATgLdGpZZZSN2kyfzTw7TFLUemrVmdwkP90IBbRl7YCHyvJESJKN
eSYd8w845dtNY1SEFwUbt9v2rd0wW68vzDaejFD11je/KMgfn50Z239WTmoBZlZJg2R726m7cxoj
ER8M4SlPAUGn1Aik/DiZk+yoqHA97wRbhADJNh70V33UxuIRyUDA3Z+yzMUoPG4Zho4ieqyTlPnR
8uHCpwxW9c6ji7BacfOMToHGHJJH+VLkMMIA/eXqnS6kKKkEUguH0FxglD7JUiXoahZAGXP4TXps
FaPmDcBuQhJ+UnrAYEqJuM7vYriLyjh7sddmROC2IV3/Mq6S+kvcRdAOOdAAOC2rJpGbDDrSeAgF
MR6TeD1cB0x8v5IMg/9U0D1iSOmyTcJPy9HNLhMZ06lMk1v3HdGdYzJQOy1LscK6wC/e3UOuWHpR
Loaxh0ttJpcGxoLF0bhlAWX8bq5X4C4M5HdsJ8mLXJY4N7o+LWjMsmTa9HTz0CNchoZjLobwsy08
mNjT4zii+rvzLkZ0p/RBcJbGM0/vMeRKasXo4hiaCtsio5MHymS/nkTkjxVPfyBUiuiUm2Glcs49
ZCMl/t+7jIq0aWhMuczm5qSBOHY1yXsriFyd6EhCdp2fTvkDVRgSeBkFxMR/LgCBNZLEPSzViMQo
3BneIrINLGem4SrhRCKBKsn7neJ+19XQzRsKMN6OmS6zxOmiA/9HE45hWdNed+IPEumPx7Dxi23S
eYKrkim1d5rmFOC2qk0NqpLD4U1KnOkXDgFuw7QGu2iUpPbsZTqjbJqMjY5QYFtp/pJljzc82u6S
UBK88kZ4nWA8SSWk5CVQ/2eihwVHpn5I/+01HBCfg4ndpLqe0nRGU4hVtk3CUmFDlHPsAnSlYwXS
WHR1+YvthlK9gHnavXn+QkCS423LsYtLWN7dpoBQyhZ0GGlFTZqYVbw/OOLcIulQTtoLq+/l/Jyx
o8+Y8A5Rf4icTHUgsj9XwzClvCU21fmf9TIpMV1Ao3Ax6OxGbZUqcifC6iSYq4Ix4OWOOSI5areH
MC/Xf02LTobH5yTUW5myldnG4zy3p+GIvWmyZ6KufLYhKPHMwiBvXpVDN0xj66+YqB7w4fCJoryS
Kex0GHs+lx9UAsfs6wbJduo8gqY8TqcV8CQrJapPKvcMRVLs/GqA8gzCTSa7Yk83Q3+kkthJb6Po
oGkbrhKrep4Iw9ewuDUjcUFhvMBcHDnOYlYa0c0dg17q2Xy1z5xNyguMrkndAlPfHm+3ZOSXcv1g
BOqR1q9nEEw81ifLwCeY3llbTrAj/6VhBPF97NSwpYZNRXhYhGVOTF05ZI1BtYJ+I5QpzdywpB/A
MuEiumyH4LlpoW32xgMyx/5cDFk+sUV+lpeYSj0UDyA1hjwoY+ItZnj+l0P7RmSE3p0yyorL8qoG
jhbSvRgxC11Ff1lpiRnbP80ySA23hmM+QOvHBFK2rAILePbE3TwHcDBMoGK38h+Nml8HLO4e2Hs3
4xGMzhhZqlEDhcLPDH9KLSjizzuNAJrNNAwnDS89ANOangyLCCn8NDvbyteOOuK1PRfX94r+RtLL
TE5/woP3/hkOgst37dkifGpGCywOSIMKEdhIOhXP2J/bu0PoXM9xpdoxm9tZHoTXDk9Bmyih1G2S
dZfwzEXhVqcSGtyH0o7R8COoVN1Nn9MJALDxxP4+xmlCGGtYtATKmOV1PXzjBt7hUBu1PSOcV8rT
0+XkCgDl62vtIcdpLsCx+SHU2wBZlvtni5VUt7Dkw9aIyr1PvcBqWNXk5ekv/Q/tUED340jFWf5m
KbuvkXlko0fjvuJek9KBtwhA+mKwnot5fGmRgFrA/qgS59fiuytEOyM4MBnZgbZGElPuR8HPw07t
QJ7kcogBQWi3K+dTNVQ83gSwl2zF45ZsSO06Esu97+bdN4SaSdAYFlxsv2dZB8fOrj1kAoez43bS
C+MUvAUurbbT69x+ILMoL2gIVdgTizY1l5808ILCGPSE8tG+zjJP3jvtEe1Zojk+OiuTlH6CQ8EJ
DFbp9n4F/kftEy1p1FV4ZEqhegcIDlvUMKUrsJN/77J2ycHaSbLAUQyc2mpY28RKm3BGoZ/ikBR7
yTnxJ3FgiLw4QH5ZRaOaa9+2OX2zmt0Eysv8AsxU7KgWGHySmm+xegyJ4I3vSgVpyLbfzkeVq+vz
8Tp64RKdkwUgVEP0+91fyTQcWoE1k88bto3vF0ebZSGRRgWaOQpviJwctt/Tow/3wv9bFSsiMLmB
HvPnDmOGVIO7DByRGEUVG6A0mZZDauOMUALvufedoEh3MecNjmnFhhpG9NIPhxC1O8RfGngEa8eP
FDIHWZPMOuuPeSKRgh0dWcpbt7A/LGktR0i54jPrVGhCy3d76PV+WB12rpZIP4gyMnUViqLtUWBZ
XAS/v3gO6ynkQ1RRrA7m8H4AWhX2Xp8cEPjGgm2N+tNKyP0Oxx+/chqVql/5KGWS0ylHQseoGlqx
UfuMj9+MSCW+3U7e+Wb/QYNMu0AFwkMAcSFXpS6v+oXz25/dGFXfJdisvaBEovhQmyKy+Af8V0C8
Ai7IkTQYyqN3/oGsQhjb8JhRrANEnU5oQLg3PZc3zIAgaXWfd3cvy74n+az+rxqhFWzZrUWzNEgK
XcXEwFpYCeZEiZ6tiIZYa7Cfw3kvHLwjt8Wo50d1mrzWcpum49atlcbFXMdIx3WuNx2pkVyY+bGo
j7t4zjwN/vrVDbz+DIXTAj9Sx8pL5aHOuRROFBZH2fXLgaySF5jsV4nYh6rxqYmFqKyRh51uQIwD
5glbeXo8cbVEh6lekml8Sj2gKM1tu5PpZ7NDbUjjxrrTGsPewv9luu7PQTisaP/FEJwudb6pnEiR
FOY9r7NNOgyUfRC8Tgc3VGsVzIjNWWf2WYteJGblwaLeRa5NUezw8GwsarUrekuHCdLHt7VN/0Gz
ZDzcpHIL8gMoNYbtSScjBNjQBP8hCax+FPpVhKyyKrx075xRhn+l+yh9mjoIn7d5MMkRCCHrX84+
wK1BxsvEeoRItl7AV19MruayRyBVKlhhF+GRGRczAtyKs6U2NEGm3oBC6QawOjdn0I2/DU9EOHIz
JpLoEvuk17A317GzORnHJ/aK4sVROMwHqD2thsMttVGaxCeqKnrrBRfQa7d7u+9Bl/mGUNP7fZK7
4ubqbdKWWYwaZZkJ4/Nt2o+gG0ajJVpsRAsgbrewUJ7xEHMzkurSs2dIt582z4Ld6WSMs7zxQOpo
1TFPaa4Dl2Yv31235VoSgcHTz8WTdBKk6t+Al8kxf7/Guue7AvAeaPl8pidFN3G8UtZ54QEnXe1K
6nh7/Sst7jOh9zurRE6qxTL96LhTt7yMBFME+46FFwk+TfMhZYFLCAIrfK5q0ryrP1+0Q3j+A2s1
YU+qe4mOhHdCO3Q71ewz+hYeShJQoq5pw28XvfkU5UY9F046HDj6jD5QBhXk73pr7DwSZAic5FPr
xBZRmEnad3TB3gDLW1ZDJaITLYZnScklMRyMbZYbaT4R8f3Go/5xLyxMIQxino5c/H8hZy1itMov
PiJesOaTu+bT9vm7kYqyVyfZS+2USxgTsgodhy697csgApGMu9IWimV7tGbQz7/FbZIhkmdh/evc
aDiysppn7aitQllFrTJUCb79iWUYptdqg7g9uJa5oMnBEj588muXl45B3sf5ZVscVi7hq1w0mDdO
vlMGZ/r3Csa4+H/W8ORZkZccPb4GFiIrRGbzO21cueucbcc5kDFjQHBG0Ld3smAZkhHcW0o3/xx/
YoNMeazcLP/tOSsqcS3SJUQQhjfnt7K32+A2TPckCMsSu5dpxhNFO62YaxiL4UzT98Iwg2DE+lRl
tS8BD7Q/D3Sv9zftHYW+xLTUjXAZ2chcvmmYQk+xQOs3g0vf1SlD6jF5LbKN2/b6fn4mKxjxSzvG
k4DnnPDdxACRZTg5+W8ZBdnipQpy2hIvCIgDStotSFpvfFsM1NjpweBG17nendc6C8MN2XJh+Que
pN1yCJRAaGNlSw5fuz1aHAIsTqIx9fgS3J9oiKG7SgAJ/J3/Og3bL1uRquFooaimldQOtM1eyfG1
hMaG7Ff/u4VhtWgF1b8igy55lBw+dZf3p5VRDI7YUEZ7L/sGlDeDjQtWjF0u2MhbyqX5PuIH19L6
OQfMeJbPEy7r9JxJnmqhs/GeDbNdBmu/ASGl4KsgIF+NWrEgtEFMhhgQ7BxXngIrBvgw4LQsm36M
Gq8InDqWVF8XrQsqeCFlpcNEbV3UTMz3bmR9ycJPiPNm4RfJCcqxHRYHPue3ua281A305xmEu4PQ
LLMD8PzP/tSjV9xiNU/tLV6puGfeEACmHWjYHL+WW5vByJCRlxIBJ7leYjTdTPTYLd9cyD5q/jYq
2881Ql/l0j90tuUqnjSyZQBaHAsvo7hYhTQflVoGfxnxkI5fD3W6T+bazieN1DDUHBjUYIn0m6vz
NgwItMJoP+pJ6sHXJBzS2+9WorC+anUSt7XtebA+Y5T+XtEg2OSj7a+EDIYiVTEkSHSpFW/HE6Ij
x3n1/RuBrQOHNuXC43xIsc0SUHsBrYfPs3EUMjqYfpZxDS1h7uM3NoNZTD0v8yKWcseoObzxUyON
ioowRYAGqMtrDuI6h57uK5+opGdSzjNRYh16VY+kRo9Xwe/Gdm+/Ie0SvsheupBm5VGBuRkm0g1X
kz/IORCoKQrn/AgM1G8mig1uuo+sC20MxejNq4zCWsuChP658h7fR7kImSH3Mo5r2gzBORqzLCLH
2F0mzdqYKLyxeyt/DrX7PIB4UJ4Go7HxILDCeHxB2q0ajWMveMXUHflnO+VvsqbE6uHUWM3MrrXH
G+RhVvGelHYYi4t5HLuuE0GvmsxFXj58DAKMp8cfQgaOuLO9MhvtelUPCVSWXOtVfq+KVq9GAPAt
fNZjo7nzd7fAoh3cwpfYXJGqFvwBo3X59JffZY87cVl2hIJE/wH/mXG7oMFUC4s8a+BqK7VfQvkb
KGJE3iSsCKl8YISeklEFhfrfWtqTDRBfQApNa+273iCKX5SRtbRPARQzLi2cmOCpCSc/bSORHnpl
2kHiantlNVvppYSOoV7d39NrG9jaJcJ8If7QXLHlGp60D6e51yakRMkx2Hx+l7iJL+0d2gISCjAJ
+gQBsc+ozM0ogs4WkdGJkJzieVc7ZddoSd81yMC5EQ18heqOmXpYp1eDEHrVyeEqTPGk/ETCPye2
FaDY/itk2HiZHhoYFVIqM3qpvIeWEBy1Jor1/0hRaZCvjtcsS2fNdDBqM6r9lp7bXQME/ZO6c6x5
hog69GFtcRM869ClgUYCjQHTuVltJCeZj1kWCqpJSr3r9CnBaHbOYaWtmGz22Sba9A6wKAuf8w1H
MUyKWilchuzE3lwucJsIOZG6cUSmV8F7JcQzvYSMH4MAuA8BlA3J7GNH5+3GVigDNFwRaf4sjUR5
iGQ4u5PLrqtzMBfjkuomZ9vu8QnSouHlghhWDwmZAVsZMixaTP3JRo63oNMnM3zRK86M+svsocQE
UGQjP7eZEpghGoYerB64j8JmW/fS7sz8XhZyJYIa3ybU2L+z9ANx02VRBk1LTj4ogvaRNGjS5pxT
MuRkgEK9SBDOID0phGCFSPVaoX5RVi8KA615TTIstW+u1qGv7gezTMn6e/4vrK7e8WKT8begNeaR
8Ve6xnXOCXEAjECMUouvniZHjXxh08/9zw589jE+k1/WVtK6KrdZyNN049xQY1yls2Gi4pPSFalM
Y6FDWnPqswYy8nj24Lii8ow2xfQKivDZKucKx/cO2Fuxq78p9kX4jyINDAt9QkcmihVIvSVEAkzg
K8IX8eOdE7mNDguzPgRrmo3Dej/RThBKLx5YkZsci8sDvePDfuT3c/7UG/2v+OiddY2w0WoWzNUY
Rd+7EAqdfFIxQRWE9PJ6NbOmMsKExpJhUySd8Q0iuHtYH7gqb96K5L5g1HUU338U29Uv6cwNBPM5
GLDNJ935AnJRZO/1UFMM2QkXZvVjuir+9HzKJJyc8/MaljLdwS32kxOCxcNyvhZxRCoy0dL2cLu+
VyABnKAKROXIYnRPyUZLaXWwVVTFMqjeo2D48ibOTx7nicPjSHRdIv7bP0l7yJEF6VxAMMBjdLJW
ufVY9j2uNq0RQa2wjw6+a+DFNlXBXBthVXP3QDASKQU1/a4BzkaWHDhWzziDZCJ0Oisq6l3sldzo
o79NQJioOVOIfjEElE+Is0nlQFz6p+Swfudkj5/wOYbE7DczOWaDGL5qE+xau/qxJ3Vw01gXC8vC
z5qBm5T6xuJRPYAzyHyJRZmR2jha3rJFb+FOXrbb90MernZOqu3ZQ00joZDsWfjDJeEQtLD0+Mmm
lQebbJjqGN3OOGmHBg8Sj0n/kSLfELgKS4V897sDOIB8gBU4HMk/+fTieK5O2EJWjVw1sTnER0pl
pEziNRTuV2cUwgxjkX7SdiU6OXdJvD2HhI0c9FBSH7at+oxBMk06A3cRPY29bCGiJ8abjzI6wf0p
ng7RiXb+bf3RvhD04E3v8f+oZJvmPpdPR0BF3A5IDQjgGbyAuMNn7jGYBAJXjrLt+K5G5TchZNW/
fJkkaFzxCZ7f8bboMESJgJ/D3Vd90d8nj50cI9QefCJ3uOmYOr4lpog4ihTseEY3S0WD1AshcRkP
VssIGWNZQ5XuraXcEqVtjWgRMK9jJe9frqNXuS3XKuxNOHltxZ8l7cUO8c+e+ADG/icy6QOjjDLQ
RxsCl4/HRjKgyNLL+lR+tvMduup11JfTpUZ08mYv78AGA0o6m1eOtR/0DuUG9jqcKKUJ5pHhdXOz
V+YIAgf6Fy208l7L194gVWVvSNCzQtAzfm+LZDCA5QnIr4UiOpSb8wCc8WEzW4pZmm70dLYFWb6v
wi6/PCvq2b4mMS2KHIlIqSlLfFnSNbk2DTDyrJQR4M75prllAwB8UXRHa6Hj6gaoaIASeoo+bow6
H08TX8bByfe5qzHZ6+mr41xrCI7sI0ulCLbul+ivireKI0StIXB1uKsWoThR7WvVd5wbboRWIWAy
rD2t8Ev/XXqIOG8wvm/C9K4NY8LoYKzMEo50gwR4GdRL4RSZD4NFKJ87NLTezbEC83+d88DQ5Mah
TsgA7M06o5FbTclrZU+mhoQGP5WXB/A241xQ40XKAQ5FRsvkM+qiZhVHFek3uNboeMILJVApUsuh
sgw4sS1y7slRPqG08gZipuBMGprXFYZLN4VRgxgOieC8A1mhkxm8hb8ELGu6aRjQ9MGkqdTfnXtI
VxbLmo520SK8r7aUrbeoOr2ETgRmOTHikFkR/KbeP/jCyYwwkYEovck45NMTujQcFqSN4YzBA2GD
vK6iba6AJSGRu+qjIRr1nu2NGfcIDis85qE6ndTAbfazNuQcV0dd0FokwAH4wC7E3KINi2lePvUX
j7egHzhxOwu9xG8BHOMu7/n66t5QaZDD/T2qB0ujGqhCuFjCFhS9PLbbCWCr5mXY8emIHhnDLrna
M+VOFRL21zGcvGjUUuncAqdm8yfC2Yglk/YaSXHye+EAV0B5BD0hP1LQu2YnBBn2UyzRjDmtC7TQ
w71yOW9TRl1VSJo2vrXO4BZp09z8EvMZ2dRCIFdCUI0jUkuYKOzmAXExRUzv+TS7xW6KQh9Vob8F
lJzJpfr/GOvMi7Xu2SSNfM13RzFRdPju9FB8SbkgiMJB6+zhVLVxC+bmxF2pFzXk7x3ZcNWR1vgG
sPPYg9JmMUIFP/56HqzkJBhGyxp9r2sGo9YeFjx4o5Zr8JS2Tcl80xn2wysndv6HNHUKA4gAKrGj
CwDftZSUkfHEbB6In+WW40LupBjfoYwLz03NIGDPpNDKNA5PDLwfBpsjwPrWfwHO1AU7rL5fa86W
2loTB7aLE0Kco8nSNBba/m3N3aJ7oYSu8I2cjFbJ23STgue+oWuhdET6Fi924aooHJji1Y5BDsZ9
o53bZ5NYGvBJufnhbxNc/bvPerIILpZbKCgPh1mvvXqODzAUxZtBf/ma9JcGhLBtMgze5uGyIsEG
GjHG2u/Q3uqj6dJc3I7vzQRa/bs1jy92UijmzK1z7C4MwjHqfXC24bY5F65td5s8yCu5U1rqJYkP
Tj9cwu3/cw07ApuouIuz5cmTGwLxjQlpykLqeiitk4X5d4LGIS3Mhy4A4HMR/z71bRSyK1x98qXr
XzlElbaiVTZwkicMutqHJ2964TzTUtoWThgqSSywKdDMwP+ECYTAxB72EEq4H9G73Crv3e2i+sqC
HkT2/s2msd5gSP3rGbmd7qtpvj6BNC5A+Abp43+LDQiKT5xVfKGxOvJ2uh/92DLPg3Uhbxh6GYgK
oIWo3cfUJkoRMICgL8YjbjrZQdbJYEk/IzN8FURVs5kKvm3VTaxT2gYsWIUHJxwydK+/3waceQTt
vnu7Vhdda4O4d4qFcxDO591EOKGn/R1WB9ITCDIfdkUk11A53we/qhqoqGIPmgVHfGn6OijVw3m7
tS11+LnPzzJARYvEzvpVOHk4XZWxMaNarU6syHV29rQlmHCgHGIyUeWCCNcOiLflAPDkimI5aO5e
PJ6Qh0+hmRa/Mzg6jYcqIETrCA9oCUS+91gk95GN4T/+/oTL86MwUJdhwpd38xkxz1CrCr5kpk7k
ARVeOUx97CPG/HU2eX2BSV/tL9wwjMxsEJGZNeulEKyP6ntczL24ER/EC7lzy1FzJRGRGAPrIatS
8COQuZhktyAjCTNquMmcYkRM/n7KfUC+nWZa89P3qPl5Nf4XK1oEPe99hZTL96hWMiG9F0mrlmBg
M1GLnWdHYBrUy/N2yxyijIYyDjp2EKT/OOBYMZUNVIQgFxne0nH9KyQlATNBQdHoxPt9VPY/005C
DOXbJZuIJtPpSkAVDGnzddlIQXXdgH761J6z+D5FQQb3Z4GIcfKAlQERPBpY4ewlVfWVaanZtGHZ
pXv6pMlhXTAWvksxnj/M7Z+Y4P1YYq5WqxhrPjPJXBaX5SyTCXBSXhVss4ekIbAGxSueOyajP/Cg
YcvMbA2TnCrn6uYJf5ivyI+enm6m+XdSh+68sL1qLTHzZCbfnziSQr8VHiHekSvYxkw/+w7EVY51
RyuAjrc7VYCdZsBWiyIKjgborNLsUjnDgSvNCPZm2Oq4fCIu++qWdutCwlc0faORux1UYysyF2P6
TUX/ypAi4apR+1ChgW39wkCK+1HAewuChovGY9YLQyoeGwvXvAbG4OimSYTIrsRNXAoXxkBXvxiY
ypDdOyTJ/8c3ntLp+jAjYOM98nISPRODJ/qw7KU5MTa94SpczB1XX15N1f1IdYH+PMorALZnErcu
QaB9PV4nrHdXYCBEy7YWYGXyaVL7NF452ibZzhpOXi0ZI1SqtqnPAsyc6ZNSPMV2au+oes+wxjf6
zbhATUvebmON9pkn1eKh4gUeMZyj3y2LcciWFLJacENK7dGFH7vG58OnBb5vFbjgZr++d3v/mGnx
ABYNErL7mRxJy6Tc7O4gOOLl+xY/RqrvaxXYOvTdYWvtZvd30ba7PeaqlxULA1WvnGn7TqIK0GT0
lM97rHNsJnx0AenJeA9xN8Y8qsPJeWYuJfh1M3xE93XQjDz/1W7w45KuGIRqlR++YuNgazrp+zqU
nMKPhlTMWJGYq2Qfm88ghLj8RIv4CBBN+0iGEOCe2e2AEqnq9P52uelKNVW8GG6QklQqxNIhI0t/
v9fhy3Qrr8bMqWTipo+k+kl/emyg1mBLq0hyW0lSBr/WDgda/7a6tUvoW19Sia6JMA0LeQH1OLrI
CKWpzsfh3WHTeUPPFYbW7UPf4Th9iqn8lI6eySqojsrdZeLoI9rm2C0uOdexTka63x4oMkoNaoiC
rAYgRcAnchuQK0uT5kj16bPFPGRs8+Y1osBiNVp7jsmzGAHuQb3+3nOQ4oaUGBrSlRO2NqHoyV9l
JZYOwD/61UV9rxLwipvR/iHcFJzUQrpiiV6vQ78OyrPbIqNdK7DtUAqYlOhdUwRaF+hVW7OpFktq
TfHkT7ag1pA4aGvuHcXiy1gtp1zlbd2GUPYfaG7y5VtviFytDJLxEnOXJw77Jg8/a39oqrA37l7B
6xo05uVk1HRB37UUIfI2g8aKhIfxQsVs94rl9E3MdvuLFrbHNzA/FgKKTcNyIUmUYMNYc9XyYqzT
Z2yszDUuWB9hc9CHwOVYbl3igcZxxwQxM7DNhxi9XziGeMx0tNf9oAOXeNJoiz1ENJs8KJOA7XxA
k9PcyvjoR3GIcc6090PRDS5MFYzja/XwOF6Vb3AbvEjMJKE+B52Qv6a4F/Zx3egRCAoMWso2PyrZ
pZRGbH7bkfuhkKuSO9H1PZUp2xhG7apta/PVM7zZs1sixmknE5CIk4HHvkrLRv1ksdOIsGBZu2cG
P6MklsoVCldKnzoI9WKLbw8t4O3VbHjOsIbkqyKIYCu/C+jVnBm6PS66GfR7Y3IoL7MBCDJpz7li
RSbJqWbCNUS1jjiGKHQrOHQjFrWL3AG1ybO2NB9fIEOG7pZ86paS67MaH5iKQ0rE96HINHT8bbWi
AaQXTMVqJvtlQJokm1xVwMerZyu1V+lgwEbSNo7SUaRYq2upr8FSGM8T4Y/OpeBdpAzrZOxGEhYD
NIH5ju+DjRZADHwYO4c8G3mN8Qbbm1mqJODM/C2yqPk54yv5qQPvZWWVQEt/pn/PYlXiYvnrmPGd
Z6JJGP8pIFe87ziFGWZxPsWvAX8mG0Dn+/SKqltkx8Zm2HFnNHHO9Pc1nhgeaWV/yxv8pgYk6X13
VJvsuzxsuPqHwHRGU96v4iZ0uD9S6K2SnbJYpe+v61O2IqjykbCzaU+6zBfyTrdkXWZjLnMGmobQ
TEnTcBLWJ9knPOwEs+Tn1eA2JQrg5JhgMce7hKXaMRTw9zMfYAWGZXBp1mWl5XolukCX5b03Tt6e
ZnJHyVtaoWg31KsOSRB2H+PHtG9AQ6HTZjT/7u+vlPBNme3Xu33KyJq0RsuyPFAGBNxhicFC0Yp1
vNWoyR1IeJWcog1ezJWmrtbLlz+TtdCWgcgRhuyvDIHzend4LPknB7myIFLMkusSN2hJGBYyKAl0
T9xahBL8Rnw561zrKmFVvBGKe7eISWoyQQ00tdkHffhDf7qaWCMNPl0HdfMhSEEzXslz5Fn6HL/o
9qgzbWwnNT4PgULPhyJBjeZ9CfVCBkHa+id1Tk3CKy7LeRLGzDc/im6bddv73l8wUSJH/dC/SbHn
Bss+gdzn3ny/RgoK2yQw0wkwnSuVbevLv9Xt/dQPihrrEfFR4D4mZz53RDxvjyQgVMdMffuk9y8w
5qbeOKK5iduRuCb3LaECykbw+LmDbrrTs6fF8NK01K9arzwg+l38Im728A8WaDY8IT8uTc3viRNP
8xeBynVgQYvG1OaDBbPwYimAGe2rWiZFgNzNU4S+vWgSTriPDoM+MYOFNhzfRG00Kr1Hk3p4wrnz
6gHk7xNhYby6/vEBuOhIqt1MPF1Aa3JzJKKXcRmMJN8Qf/x85gdPYJzxVxOL6hLUoqpf+X56Is4B
vToPatACd6FDxixITtnm0w2+k8hK965BUzX2BSOXRv5UGmo7CroEl6gbcqDw9SaDKcgB7ktIMvCI
v4L5o1rKJunJs3UdVnMG5eTTKs0H9lyY76wq12XIOrs9GoCuj2Mw3DUrcHUZHqRgH4KcsCj2RQAj
C4DcKRkuH0G69YlPc75RQ9VcSvVsn47zK9bUYnlu9o0fdKxxRAK4jC4C+6OsrgwvycMC2WxiJoiE
icOV/QnaC9vLYv4NjhqAIZ98XZvyPKGn7cQKUITuN5Ud8iwkmadd/xQ0oDrROgMui30g/9k48Pbs
ZQIQDMKj7fd0jEJuqY5ernhV+deQ6h5pzKoYrEAKExkMLc/vHaiMbeKrdv1ZgBj14h3NNZmxvzUv
f/o2O3bb5khFookwWHYfiNg/9M6GkxtDkxD7u4NFtK6Nwv5+GHPnYn5IzKqtV5s81s1QWbRfd6aq
II3bqjunK4Yfl7lF7WKi149mL+K7GOcAwbwXqXKngGmrnS4ItLi5UdsNHlPtxAuRJBVIpljsczuo
nPTrdHLq64t/PBFs8UNcozpStmhBTHBNgLRE/yfnC2UShfcp+DUllH9bmswHQ6xLuiKIP/Eos32L
A3OndpjpSWL3pPCGflWPoYHnZJxH+VgzqhZudR3/spzsmBLlBQJ2J8uhTUS/Guj+/RvAQhaZkD5m
qnBXziVZIb0qtya8O25g49ZMId2rP67HCtulI88jgl+dJHVm599EDybMb0vSvzyuTOwAr5+IZmWB
vlXcyTnvdkv4maVnJ+k4DrLsL9cFfIeRoRy7pKFvKDXvaHiBK87zGZiQ+k5ejcRWzAODPIhoCOB3
vrlLzmAcMaOx6ExIgH4A4o896gYQEZn5GyeoIcJLNhFudHhz38yMZzSVfi8et1oHpoUaOqS0VviD
hoWPfZP1t6nag8IfXFeGfvyBA0I/E6HPVmCapw9fTF3DMC/SXK/B+ilYM8L5BHyotYx43fNphRBj
WjzDcaEES4eMH/mT55/eYaYUwvsQA/uwoB1QjcjWRcJp76Igjqcb7aWWySB8pos60hhMQLCai7Ho
KM/IgEIKfOeWAfgzaQNq7TdNYvDQ++sc6qD/wWq3no5FwWYbJYbvqIuCzby3eHtHvT4tEyuec4qj
APy8TOzB/zVIftZThhNNunjlN3q86XQ0yjIZVh13m13ZZUNo76rOD6BNZzcf157c3khfaOe5DkiU
05jAL9VK1JpxMz2heBNNGyEMN6ZCcorcadKh0XHa3taRETdOXjcB54Wzt9rVG0MCqkbYfTttHB38
9vUOKrcBZAdhKPRzCfusx7ZHhOd1DCUErlAD9B1ARS+XpDj151DoenxAf3h2UNWaPs/4z22jJAfT
tGOFHgI7nZTg/OZMJmXZNLFkZmoDqEzANxH8pGzjvqXnI1y11mc/SEDZ8lNfNeVhqN5rK9gS4F/H
SHtIkLRMXwJCC0NCsG5dSRbdEFypri19xTgc3MFyaRijEFe6Y4h6BYRicBEZ6rYdSX+KQO6FyO2U
/HGVHJyHmr8nOMzp9/GsFywvIOLwGZngv0HWCh6dxSPKkf0ITwnIQKfmqcep/y/ZYl0iG7IpQkdY
Du8Xyy3DMhK4XEN//7pA0E2hFHJAtjMeDGNhoIFBZDOvrI2ABY1AJeadxUP1iJbbc/fXz9ZXi/xy
N4JU2VXDSbv3aQWYqSDMp8+YFWkYkQEDFvzx+2+ZIkgGcqUY2BTwT2EbEru/VHb88+7oEClyy8dz
o0E5sxJ2B1rNess2rnsBZbNOe9yQq4+q4Ena4xjGPsplLcLQMY0ERvF4bmeCy/Nv1lZTdlms1zzR
HgTlgLqbFkJgk6zILDbeWzvqNQYkFeERGiXymtsXPNcMLZPwhkxrjO7/+Ivurh2tqy1qFFKLQyr9
29geBpHZaTo2zfkixLGbtSpz7t2Xlo2WQio3EP2AebbtDb02+C+Vx0rMPSkgpIT8vkITlYe12tE0
3klHxoKs2vyVL/4sqUaHgUCYag10/Zg0tA7/yeRd2NAVtqvQTKlUXl4uj2cpWk+Mpk2UjmLWRaHe
PWdqHFaxVXUjUG7Yv4zKiNW72eDx8YPrTQXGYtGJTWFosh9zeFm24uv5U/e4WXwu9wajOyBatk3H
XevYf+pZa0y2wfvYC0RzOIFLVrh9h88PaTWR924UEcUrqKgZrfDmiwGtiH423TZgfpLSPeG8EiYS
KYnY2/+NKDCFaObyrsQjm2Y5nDSDavSoqC9LxhpOwoWH1gfSBos4F1su1QicJMBQcf+6GJfnSusU
YA3gSuCuArhpG3RGF0amfnjfACRzZXVGPxCsBL2qv4oJELf1GIgYgBAMVF9663Nau4FNIoVEi3u5
l6f2cSCrfk6NogNOHT0bbVpp/DqeRvz8N77zp2o96DG5pH1TBDYIuD3b8KIuSTuim1lqrxWgwbo3
4p9RT2jaG6tIjRe4M16oo4IrlF7equlyNHt9EDOi5NIHVXK5NuO7F6JQlpLd/LVDuFxFC0PbtRby
rTn84ObAL5g5ZW3DqqP0j+oGDf1k5q0AdAZr0n6M/zocS/g9IipUrdMZsop6Gx6mVNp1SWAIts1M
XzuAQbD8Z3ZR99pgpk3xwU3ATygC6G/6zPd/Qxro+sXUxUXVnbujqMW8iKpaSGO1+xtN0lnM/PIy
uj3xwbvY+TXegg5S2XKCCSaCCZHp2ISZtusLSK7q2WFBeO8JNbykp5Mvmdc6fMvVt75fMA553iOb
EWMm08xX9kyF9Ivyz10pJRfshzLOgydKbLuTfP73grxICJSu1BAeWYGXXOMchD7CPyfUM6FCgrtz
sZkV7PfYsfRYqWkLBR9PXP+TCv4htHpCp7Waa2e9tI/EL6aJffW9z5qSqfvoggjYG9XKbfXdVetg
3HEfERntumBaFK+e9rKWRadUr0YADptMkJw5rJLD1q92qd5Kr9LC/J/HosJCzBKVxqYuVFBDhEXu
i/gaXDNbfJSZRt4PfTdLZtZNLrp0BuYTgEe2HM4ShWrB5tRIbRY64alEZn3cpv+cEe1Q3mySwgSA
z+1cD4nHHB7hexzV8tZAf3GYa2iQgd06coRuDz9Mork0rdPP6pliv7HvIG4Qh2ehPDdLSWDHEpPl
klZlml8sYgztyN4Stz/YkXySKTjmWwgbC6y2emsxO5YMt3ZWU+exDRXOyzFf1wl6y9+iHcnI7BJA
FoZ8T4iJkQts1JpkLaPTtmvrPc+Xvi7yDmBF6r2E9QuCiq4r4KZf5Qa+iqJLBqSSsHqV49vFsey2
O2nCzIJB51vWTdfJeqrbwtWQA6Y3YoeeXubBLZq53vGRwzUBvLyyFw1H9pjNgY937vHAk1c00LEZ
mjrnFg6Y2gqMiRdB8A1i6CThoiMRT4/tXk9/ed85Xh0Mz0ESNE0oAiKoHMBdF3fcqxPdAYIwwqQ2
TnNvYwwX4pmqoKG44rzKPYJBRXLs4O0s1Hgh6geESnUrzX+NyPPpQd2JnIKd3KTb1zTJYZCzYFJZ
wFpfCTpwlCycVsJcdbxg0TSjdNoTJrcD6EAO5sz0Ku1l0VH47bSgD+6+2FiVavBCd8qFy/f2Qrp+
LNGTYpCizen3qKLeau4kb2Vhe59Bz8xBuDD+P2D/b2abldGN9n8m/bN20QZ6RdauUreZpFDdrQeS
Z811aXHByE0SuHMqoLgq989YGLzi7SqHTY6U8CH+6FSZBlFhS1+VAm4k0E7qQbnl6uDHy3sZ7GgZ
RWc6l62rnhk8hR/xmaStee9+Oi2tbMQnZ3l30NlMxAaQOPVJzH8tsqWaLKnGojivX5234FJJ6QSs
yRhDzDORTYpPU5PYl2oknxZ1Mh7oDYEHaOcNKl5AVHdgYQOqo3YKfrfopotVLWMUEegAJ6oR4yd1
0WA39hevpLTsinXlG6cCdEpVZAJfEfTaL+vdyhTVoZTNPUhcOYBUbpwyrD2zaUIP2IKwJBjJgqOm
0NfO/u5H7DPxKR/M+ly9RjA0RizU0PJNIj5UEwhW59GCFlhXAkvmaZMLVIFRroR9YHy/UjKDfArc
NGXnWokAG+ogaHisF1ONxkPlFADkQ8ys3N5neiZw1VhU6KZT3nKVBxLL0xbZFWfHKhG77b4BlUqc
pmZIEKJUHYNbP1T4Ax1NtPZUZm2OVxLVoTP/+1Jl4q6WG8zYIgnmnAgBEFtl7fdbDdy9yI9/aD7a
bieVFy3hcXJ+uCTmTP1ztC88E1+ETyiwKGDDU9R/UwPqN39ALamPiFD8BKbPa09Ei3S8YIvNyTkA
I1ZbvseoTUbYMvoEDjcX7mFAQKK2WoaTjO2aN1L7J58N18ZSFBTJfXBVme9EA8zwzFO2bTK7kGLK
u38cvkzDMyGrgLaeom9MkBIq1CVMH1QewBFMHw4zlTLplnnJ4mr8sX24t/UsORmQMNEjIPywECJ+
uxZhlea4h2AyYGh2ptzYXSCrct3S882MLpQAd8Qe7NC9WXKsHcWLV8GOljImWjHjfmSLIThfrLCP
uEe768b4ZGiUNtVyNEDJ+FVI7ea/2tJ7goad/wcNAFkNie4LXyoqpSsjatNbfcxdxHOxFRxlbAa8
c15QpE1U45/OTabuX7RE2b4wYA/cZG/YtAB2Pdl012WED5xSPGK8laZOEfQXOj/iI4Svga+Uk8yp
Asg+6mwjePWNahRZV/cGqMpFm6GVQCDdXIDCVZBiHLvUBWmr8qV0zEi10EzbL/dXg2V2ZmTsD/0u
UmNHUzjy79N7r2rp74wFA/OQO/HtwUVXFd1/aZDa/0JOR6STG4Z/OyH0tyLLcIMSJt9Rgg5L0nWq
GKiSWN+l8dYshqYgnxTSBNeyBcFggAU93pXD9sy16X5Kg4pARBjq4VUSnZhQQgaX7rURe3RStyAt
05TIZdzbYtyUL0XD0oQsKE1OYVQW6atMlMNNjBGYpP9vIC3jQjBx30K9NQsiRI94LL0scexBuI0a
xcWK/mmBX6MQVBGTsswraYzSLkLTFVNwKCii9yI4jy/qoRtK/JdWNuSpOQQIdFJe6mfMMYfJaG5Q
UoDZbuEYNFd/r7g6b5rst0d9nl0NPSENvAFgg/2xrS+8xTx/KCyf9UALvG3sjpZ58V+Yg9KghA7M
6fuzQ8HP96dccNhcfdXe1IU9CX5OfFOfXpzXeppsr4wQakhZ/DKim0huduMO12qE7f2UaQ3UOXCM
QobbpwHckpPOap1C2+RHEwqyTiiw2NuyLg4oXkYRL/3pVZeMcIBLZp9aHBzZag4GMhwTEdsN1KEd
88BkUYEVzJqSP54tEABqT3HkFHofXXhCP+KUYEaUSYzMSu6jqwfbprM75b4wHe5gqmFZskrupVHn
KI5ObZTCn5aYrSCR3eojTKA1aqK/vUy4h0jMvVo9MTncXnKIDCYWBjbD2nYcfmDVCvA5vFcubo5a
2eGxalXuPdDR6kch+vdWwF0mxx5ib1hphWcL5pP2xz0hhKA7yAxgeu9/BOAdFhOkpwIBXCrV5XYT
PsZbF/smK1pHCZmshvsnDuASbw+9SlvI6C4vwbn0nvMwuCXvW6GTjmEHeNeEsoF9WZNvqCiloarX
UA46mXGCB8tkkJe7nX9UaaCjcGUNNCCM5ElAjjMN2x4LmhkxrcpekQ++jHhz3PYEn0BqBTKECgwc
tIYHI8t8dZjdyAdXY0Tvz4W1W7yrT4wpooG/vu+SgStBMvA0JuDEr6jdU9LYqbvmV/AAOXQJ1sO1
Ncr/ihhWcmAadVxylo3WOkfNGLCUTrGzr/+1ZFRTi6h+1VNxQcxBF2R1Ndu+Bf25aBRcoMmvrRPJ
xzCbtOUpcLFE3dFTEk20GeH88kLySkkJDcLyzOsoDl0cpVILR6oDBHnDt7VhrftfropObeghUMGT
1+bar4iV+ijky13X0FMcGJSkis7rYRTvMvb12TYMpAhAiUOKD4c0zWVwDucaqthSNcvsekUZaFbF
ZMLsrFCQk5mMT8xumq1wInrnwSLOMxvrvpSRC2PRsGSnoLmXGEafoGMRNIHV7g4AjcOQdHbiWKPL
eYR72yxNpj11fkJC+nXGybVMyJ5ePHDtb5O5hPUyEMyoQx7rwNNkTIP1myANA2SS/k7JLo93gSH6
vKSmoiEEljKQsjoLxEKTTaPA+UWQwo0BbVASzcFgk5K1fNkltyt4vX2clxNrQHg8UdLP4mPHC3+3
/U/Cd6Ses77/lAzRnS5Rj+aEQIX9QNBCfZDHPCKcV2QVcwXc2p8lFDPVaxnz9oDXfqhYx/uc2SN7
6RbQmGe2CDB3Y4d4bDODBbIC2ClcdjsCCRMRXUeXO/FsvjI2vSU9m5jojyHp0P5Wxfbg1RLhXQOA
1bLRiTym/IqBCYYZ6V6Trbqr5YSHjW/OVLTDcjt25m5eA4DfKZJlbFVFLa51uTVskrLigZF+yI3w
9cZRR9YX+iN/G9y1SHtFANmg/JVX5P/ZmMduOT8c8JAm7kfQqWzSh8O+gUxpqU6n0xZ0A0VhKuYC
kV1s4D0Vvohd96ed1hOZ4r4/fg1lbytW5VI+wyEEDkkKsMdED38YvBlOag77sX+Aj6879RA6n2VW
Xi2cXlJ3dU90UCk6wl7TbOdS+CIM0SrbVxIyvY39UCjpuTO//8GagENwu24QUjlEfCv+lFqSPkVI
yfal06C8D+RmuhcTUJ2vF3smEafHIdaqJgdkj+5A9FdA5hUKAbgMWPQqYNB/i+/C6vxpjftGaBL/
2md+/85y0aCCG9dHyPLG71TkhV3lAS5lGDcU6pRlz8vb2D4eTjoXDRZH+f1aN9ZJvJzZ+U0Gs1Yv
6hTRO5OI/SFH+WO8OKzVHh/WrBWuEyKvsDqpHpWOhk6cPChaha20hE4b29jxLspL5Rr9UBkvVfjk
dzb001BNv6dLSL/dgx/SXBbqUevmHl1AY088rQFUiyRol/uc3jv6dJyd5avHXkD7PIxZ7rRZAGq/
o4WeNiF7qIG1Up5/pRue6W3F6H9575BHju8pYMKUtSuDcT0jIF/ShZumQ0pkUICxK96isH6ziCI6
r5DV504nCvvR5nXZjZqHoED7xrrbEGBKcuesPtvE3UHDBPecigHsM3zi/p7rOR9k5ejDejQ/an9A
NPBClUE91JuWKT9GfDa4/Vq/41crD1Y7INodjj8lpE5pAPANzftZvr9twnh7NE0VnR+1acJDFhCy
tlw49m1TKgN7gaubTkj5B3pCj6PyXpmH3wtlHbi/DyyV8z2B3j5MEoBYibbVPeC2aleBVd+1WXw9
09lymWp0IKQiSZdB7KmogM7g0MsEFiXZHmNVPMeDhbl4YobXJXh1B4ncqldRG85bz0e+POEND1Bc
rI5cvc2IubnaU6zqpkaWNVYZ/b4K9IHSgwDutH/0QKLBNYTWliYZziXive0nnsspDlZZRqp57G3g
LZrrOCuTpe1SaEtbLigIPbsOzNodNs+8Um407CH0PmjRxUPxMv0nDaKxb/Jo2VfIU2leuIhxwVHN
W/72955Qbrr7Keyv+ZAI/KTCSugwkaRGCtUss7cH+65pBwebewqfLpu9Mckr58Xzhwqsx0kHGCKV
PwrXgaGznsau/0BQzmrNsGA5jcXLrn3V0RROOdEebwzLwZ5b3yLOiqkWu+Igimg/eN8XySq6gnXO
X+KGkYrxFg1wIMF+5eamNYibyS3V2H9HCl3V3UiIgpQuY+yWoyWkd0xxp9EjYXyYavU2jWHx5Y2i
f319xO91bILuMqiGxlUgzVfQX2gtVCjcGjMUhtpwyJ6J3HdT/R0CMvos5S456vvKqFVNqvWFjCpb
YrCbhclWpHZivCKi4gXqr+Vzgf9uhLlJgHv5QSAKNsrUKQns4IVLmrH/k0k3+58sxdPmBnyeBHMv
EedkzSPkPEYbz2qVc40YIuIehmnz66rzOJnBnvoW+xPoyK8R1kkt2i/93mU3gdgR0b8/8ZrDXcP1
1KKR7Ac5p8cHPbM7oox/oltYP+wMoExD+ExISDe4EN6H6ektMGvF2R96OYsCa4ZpU0Aum5wg9rBu
+BuZDHXpEJX5O53/PEd3uKAlsExakUYEybTEQUFzWttEaMGXUUAopMyYgJf9LBTi+OeBTSF373BX
mo7ij/a3CmL//cGj5nynNk/hC+K8RCEUTPcp1mv7TT0uR9hDtwAgHklVfr+ZTXsgm01IPItSFKxd
kQAZEzyqchzRHK7Glx7QP+3ufHBoA52FRGK50aa9OCBqdNIW8n8Oe0sltsPCyryjn0YnW9ryqgsz
EdICt5f9nj2jdnGdERIeLUYhsRX9swHz7A3weR5Wh+M4oM5bFRfRNhzOoCifpEKPYvwXJ0PQhIGp
J164KIg83SlSyyMKBqcBBXyY177JzCZL1oqedr6MouRpUGRArl19Uw1kOOu435L9g6LCKK3lyojj
jj/Mc6B2+i+VW9tQppwvd9gGGly6VG/bSmH12FYoNkIWZNQXa0DBRI02+J6usu5f+ovTzqszP8cu
PrlsX8wW25RovEaQhfXTqF4/o7J1qcm+Zi81EAMdKtcEV31v71q348A8GBMOfoOgASXWer6lOxcE
F7GX+5j5yrMIM+CvjyT7WfCmRfgzOD/bMswFMawzXWqvKQf1NMTGQqkxseiTBrWPrGidqrAnxO2Q
OmIE7FnJ8Ldi6Is3O25sP23KUaBw8GpY6GfieAZm2GnL25UH/fg33pCNGE/YZizFNSTpLE4ZcxVR
lt0d8Z28GXztDWPRAzpynxODHKTGSdqty2+B//RRpchj1nI30Bp3SneRbcz3bsjJxVLln+/+hFQ5
hCKxJnHIPNCN3Zxwc7T2E2IDM3ine7NzDleRi0LhO7CH25bGBB8UDPz4o4/8dcf8mDrjISZXamgG
I0sX3IJEijZ9D4RwK/TGKMywW7lRRi4GyR/BUs+IzuTjC6Mx9Pgl5Y1h9mHgknPJYecCU9qzM6nt
D3rNvhXeoF15hm57MQ6KSX4e54N7CcuYoeM4EzbCWNi+vcb2PHqiNCmthNJ23XfSkIdzDyp6qlen
d7eYfui4syepCWqKxwMhxSjeAsDlxPdtnHVYpr7esouieGLQA3i3S3UQD/VbcOi/2r0POv6leWuU
DaOoNdvPHuvSLoacFkpnLdV1EEtPUhFdIymPYAmtORfY0QrjhqF2CsVkXdJs2ZidKrMuyePIxfNr
04FQfU9c0fPRsWyKOKZuouDiMV3Ox38lGAVoVS0B1OTCS/iYofRmQbs6UXos6a8gEJpuwa/KWuXX
r+TT1u7skqTuO69ggQljGHn8HL5HpXfXEsJTjuM949E8WLWg7QAQ4gDkh7QVMutY6UoOnu3Lreju
3n4+I87V+PNEkJA3OafWr3fbbyIKUWmMfkaDOrEHpzuoIqSPJTk7aPAJc3pM02TcDufOuM3jpKcU
hyHZ+OObCHCtbbkimJKfx3hNyj3PlViFmNQOZG15rTmF8kSweF/j92qY6DC3lbg/p8keY4pOzXge
mdOPrLssZeNOxo2hgqbkpVZ0mnPoXN5Br05nXgUg3qUbTAqcdiB/SztL5BCXgDV3zOg83JFD7Nd6
dqiGp1nT4mSiYfLhDj9Z9O60pO3dHR/YyT+GHMs5pHM1H3DibhBPDYOJWex9wCPITzW8ePJ1wtP5
13WaxApPJleMVYNIHgD9cpyKbuiDHAby3jP6y8AhzBFSf1jJ5JFskXkQX3vYG8Erd0/gJVcaP/9D
/GesqcU4Q/bx/DM7VtPS78tYbo4O43HmRK9njdzv2UQS27wc1YlPySesvfLAIS0QlJXOAVUkJIYa
6fMn2Srh+oQD/xIA5iwHuKPzwnJ1xoAdihYQE8fEeyANriwxyKw/Z0ZDtGst2lwAj+1doW8uzKBy
vPVai8TLqCIieIlMCepo3aaB4AHAfhqu23JOVyIEejt0ib4rDsU59UxdV9UEZE54dWWVeFfEVFXB
lm4vUGdIav/iXDpmjzgNsy4AQkgS01gHHlvAmdXV4gwPK2zAv7rhO5ibPaTss5eY+cnVP2dAxPvQ
FFKt3pZq1/9fgkhhdlbJBOpr53G5Zq9//7vqMlbFxvQ++XT/fgXZXyr4MLKGA7+RApzpriyFZnnj
wNCXeI9RtM/AUpHIxs1srHXqa/CKt99IKSumcFssEiiftTVatlPQMXLg+FqKjwzXW4y5SCrWr9e5
IE4Qipu5hGMv/BKW2X1tuRBxA8x7SRyoOyFgoNSpM9+eMqQN5FQv0VQtwxUffNUN21PnJu5PQH79
1TLYfSaNnWwhyNZsUP4xUyPocqDg3ci6G31cmFVcU6TbIk1UdmPmNa2GTpDoe1oYpUwRvJfYdMX1
rmUzPwCrPpZbqsiYILPFl/HQsenPmik0unVruTIRnqG6snckkbrWxG8CQ4/Aq+tEsANrUntkoXHl
S6DYZPtW4/1qjbH+O0WF+EeioaQhDMvjFBY17FfcDaDSIwXmfDdrY564plzGqRwH1Ns3JrnB3D5Y
YbeEHyfW7jD0XDoJBrHr4xsES1/AvQ2HfSVTjc7x6+h2PJrqrnJAdbK6CLYoLoYxLJJLqBGvO9es
82ClpC9pRC94c+NSW8FSy8zVpCY+VVXrNuP8NbPE5uYQme6ZscQqpo/sstLxI+dB5YI9XwNGROSz
It8T+phnc0ustzcxCdQlLxV7SkFtQKqO0YJJbZXSnFXQATMU5ShoSMj0DiTc0KEl4m7z7oQNiqec
B/rXAGUSvG9zJ4ijYZUgL9pn8GzNv9V3VWGqvJt+u0x5zLZBAtxnV+GD5WvVPcM49SW83x1wMla7
E9JQ6afRH7RmioHac6w2EnnRKwzUuncIGy3Ej27TzPgA6zicJMD3kSOxu/SgHJOb8oguacJUMwLc
DyO4Y25CA+y/cBFbIgoUr9p5UWhjVZ7JQUj9oyfrUwu7AkMnD1noLNPwTnjKmvjzObcC09kILGTG
TPnDPZ7aV3OhMi2LhBvN6gD+T9y/Jjvm/rqWsI69a6+1n8gJwLZso8kpvcy+ET+WCmYACMg7vJ3V
do7cZ5FfDAX+0jUOM6TgMT2W4NAM8n+TU1IkFaTc5WNq0MEeUbZUGdH+FKePsCVbEauYtJHN/hO7
Nano8DULVb/mBTqfdDFU/Cs7YCSEtj5/CaxHrzQDHrs3foVSdwVuMjjcB7yV8y9ayI2dFbsi4EMW
AoWGvVopEHYAvTVjxfM+TtaTWXFAzdMEybqPyVyZm010fKqt4LIHZJtpN1BkcawUarb7IXNflloG
ecuPqd+EWklVVaYBynFI8s+GqaNj/XHaaGBmwi3A8M2o0I0fdOfbL1HGWC2NRkPia4CzN0InhNYM
fEOsnfgdzNfS2b/zhrSwRh/eg5M4bi2M9dN8W2xtgi2Yo028/z8BcH95g3Mj5EbOuo4lSt9LhjiF
72DIuym6fXV3HIaOW6ln52ktf6gJMNh/AC1gGLzfVoxohOSV3BOiSz4myGy4LyUFCKQIe142mXj7
WyBn2HWCAsfsKAHU3eG0mrVudiXGEuc0tSxi+MG+C0r0PD+vwn6oTPS2zmjG9NVklsJtfNBeIX9+
RImrQtKJ8MQtVRCN5LpWQ8A/Y3VzxMROOyfkSJgs1bG5KI7MBIxYvUe+GGbSwx0QzSmVj3zqc76n
T0RvvEU7S2mmqV47ni3r0ASD4pIetj28zuP9KA8RnFzcZhNVrUbs+Y2QvhRndJ1oswRtU5PDZIDO
cH1juSV8RrabKlOGhknAZeSwJojx+C0nGRUh1G0L+QTrMaulViKoXuLjszsorZRuI15v2I62tVXP
JcGCHkL8YjanBerF2s+z8My47+by/KdsDYORFUjTVo4s5eHh3Q3rij6t8Ant+wKogdFE4HF5LqhC
Lr2kuPJnJLV6qHyTkcAUas/61rnR5H6q+FAsBaMkoi2BuUJ4d26+OK0NV06o04Gz58BQQSC/zPZJ
iWwgTeYPL/wYI+iF2W9ZowT5qOdgmmBeOTBiuAhR/XZZiP+pSbaw096DkS3u/ATqFAkVzksFf9oB
CSRESJ2u74igaFTH62GVsEsYjVJb92daDFem1QpEMlecdAeCs5MJV7ufex6d4OT16kBHNSbtfPbn
x96/++t8u77wP/O9mESHD1Q1vTHn+eyzTwla/diVy4VGwuYE5EKazU7PJsxrfNBnT7Abft+MiWoW
p/iRlmd58OHpKMuJlpil1IP9x6jkQxa3p/u0ScAAJNa3Aguw28YE4EWX8VjU9rgA6vC1/uM4Zm+n
kb5QeTxSGU8mS2fLJ+Emyv00F8mdwP7t6n7CFY1UyvZnkRa0UAavh4f5sjLF3BvkuvV8xVOgNq5p
67y4C/zoN4pZE2RpSHI7S0VlbkinGzBDUW5pjXa3RwXi4sREYvu/QVZ1R2ztDxTqFMYVRM8O0JPs
M58Nxsir4yb82u2T60vv0o4nJh+Dh8vSLCVSuV54sGKQ5tAwldCodqzUmv5Avz24lh+F4V88YV9T
8kOAObvsjsQ/I0qr06uLa41Lntgu+cgStKeRUh8OiamM82pwfkgMgUh23fNnNUwTGoo6fZDMuS81
fYM5INNFDAShBmtdUaWinG/laIHUn7/XCEWKkuinybh8omF7ncv6tAE+SmFhMrcG+4r6E4vt0AAc
PFEt53uFx3Q6+oJ9anmvXEGshNDFZVcghKj7rogVrNrfFecoKtDCPSU67D2LqG3hEk4iX6eICTIB
txcGjOZNbwpBMw+3fE68HbQjK0/g0Oh/8ESkjYtCFhq4w5Y8UDilHTFqa7ZKDNzV9qaOYI76Rk5m
KLsemhoX6h/AO1ajgVn3HIVC8Jp7J9LKNNNlKMstiUzXJx7Kla8gnml6meVcVROfVOQewV7fIQWC
bXewlyy4ZOfqfyNXD923UFACICsL+DdN+XoLVMb5YUtzdLZjtoDZnL3bddsyuFoXCc5XK8LLxaf7
LgyY/Sjpq0HVamHeFg8Z76rm+p/EAa7PKhj8gcykxfBoGxM0V0BGhpEaUNW4YzDuka4jEOsTbtzy
JKdE830g7OMvMO74Z+DA4vPnleaw2jd92ylP741yj16dbqVj/fsZ7tnEFs3v00hBT9RVQ7ViiyEN
NG1pETKp72z6wzFtzjUt8lCj3pV8z8a0KOxKbOV5qjtwC1USgu2hgJeldCB9vSasLeMliwuV6nCI
0MXLl6NphsSYfbdj3+LgizU3346A43xlAQ9z2b2d3/MVuRRbO00Hb5CWitNsGEmJjlCvoqrn7bNX
DCKKk+XoXI9YcRA/vA9OnAGhwzWttk21Jak//5d+w5BkJEsLIAflVPH453ocBjv7hvWbLkiIGcQ2
huwaTMXYgS/a/X6chEQWday0bpLVYXEZWWghihz0KFGMZ9UDYST3j1ycuWUuutDTodzWh1UdvYyE
rM9u/BBkvJEqRpgf61+haQPDtrsFowrteDnPebweewVOJZQ+I27teTC1Bb4pVtF1vvjLGG0KWR9x
CB7D5ziNAn7Roh7osXLxVLZGp/3Y8TXB/C8s/JRjJqDoQzB45AI68KF1DNBw4EYXp2RRGKwQenrX
E1cBCE7qzZboDA5RTCs6L/I9TIGbNim5swEVne1nXjqmVK1DEz7clm0nuLwg8uUF3hLS1ss+4Qcp
0axY0UsKkbXaQboJxqLAGHAjZ7ob5KKinNbTkHSICPi6pqzqG8kStlooc+WmNmfS6fKy5ZcfSWe2
qa05kUmjana4OotAZze682h/MOAVd3t1FHKM8HKdJfKfT6tqdTYr7mOT4mp5/lRSd0QMqWlvxFhL
8TfkqZ9SKyufAoccWfOerSOwIwUJKkUTn+OqbOyli/J/pKurYIPc/5O0rlp1XmvioFE7CBya9QWE
W4P4kG8CxPvlIJTtIr62KE/xR8jUheXTp+ismvi9mSsAB++HqankW12odb1tC041wJWV5+hYFT7o
MCkTxAeTW74BHemW4tFS9GsLYY+m5FtuFuv5HmkAshZjDf3wdMIjUU6uNz9qUq8aiKFcSizD8J5b
IDc5G7f+yN6NcCmBqD94BdjtrIB2THiKx+lfdNjoyPEfo6ETaSAqRW+z/wnJn1x+IAEllTSl7Sv+
1nvEnad+AatxDuF0+bQyz/n3Pz/6lXRV+zvcNYD2DQ9kYnut2pBYaa1n4yy03hWKOV/+rsul3pkN
p+WotUyYLcOxy+DHeeCkjVFhsYaM67avBuXf77RZorZat46kkGtZbonNSoPvcQ2s+IZdTTsg0oPx
Xhdx89UNedCGlFKRjjqZ90uVPkjj1BaapmknMBKmIJ5lYVr2SCQ/SkeZKzBe+c7LTN9wXu9fguA8
hwmROk7lHp0Q8lxKx8Mw25AmvIuLvpP3NivPvkKvUaFIeywM6W6osWWxNl3R78+8+1L3po32OJF1
lJ4hKo/01kMwXQLbUPHCYXl3LW11l+AGLcVWAH/P3Gv47RaMWsZ8aCoLO5TOkkDg4hhhKuzrNcU3
g6IyQGGoIhnxjdCZijWJ0bCQL0elqryumHKPLpDxAtNHB9Lfj3IFDVpNlHMRHYzJnKyXncVdgRdI
RwEIidxBV9DcISUiA88vKc1T1FMOd3m5CmkeLxYOqA3bQhbVclb1asbxcfCfES03OeKsIsiD9p/T
8HakdEZatiVM0Ha6nBV1PzMwZUfCxrX4Gyd3oV9TpEexkdr1SW3fbEBWkPe69jfd7F+53TTuSRvD
j0tgVI2ICrbyxRWr4F82H2wOA7ezfMsxIjUxFgQWMAtRtaifjyRZdbKoN4IstZypqV6iwvOwnQYK
M0SnMVSnWH1pSK4vwZB31U98dvUkiHR8E+silz6c5UN0TxW8igRv5iCvcYu0/J/hXF3F4UJ6EmeQ
nNLd2TM41Lwh2Jr9LvMaL4AllPCwm1nB/Wk/vGQ9UrrwN7Prym1FqA0L9vBPmjHSEIh04zyZOfsz
1a3ZM+g4dMYF/7hXOg3v5LYh4JnMIAp5XvBD6YdEguSQH2gSY/1tMKUQYycfEgmKPLrGZjIobMqx
vx75v6aHeiMN4vws1xUVj9TmRYr1YyJTPfsVz79bYqYOVgYtm/tO3q17yK1oOGAAYNlzb45lvUcj
M06YpBTK7laSeMVDj2v2uSMji2S9ILB5xo3Z6A8bmHU4RmLBsi0TIIi0/Bp/RkLjUqh5aCkS/0zC
NJ3vx18CAl02t+iS8Q9fCeJNtMgyUaLosBqw3zDZxCq4anN8DpbntsP35jt1hyVMtXXXHSjoQFSk
nlqGcrGZn+ne2hFnN85pLfLL2ACGohgH1Hm8+GdOwzzOOHr6L55cekuhNbVJmELt+xjTXoajcFzv
LmZaTg+/ICY+ukmS4jsRxWwmZ5sJ0A41lC4cLm7APinc19Q8JoLUr4dkLTBLhMVRsx0BwlQRi7W6
0HRfD/u5APfyTV9ZPOPLUL1tMgfLtMSN7EXwO+0cqNOsVasYeVijsiF3bVQjDFYoN9e3bMpTV+lS
O4otgxwwcmU6T4gw0eS2s53G4nSOlxhgneZgu/GI99uRlgPEpsSS71kjxogrEeNeisARpEcdicIA
0e9AkX23fm4i9HA9sF9GiwImQ4px7Q9IOjKXXHWcnTHoU2HYcWsVfZ5OoLQnmzio35FRSe2tIwHn
K4eqJ4hVEw9r7lzlcKwhRw4ymGWpD/zU2wvIjr49GrVfpEsWrrP+On0hmib71YvqCvB62DwKYkvV
JvwbnS3IgSQ4B8nGEnkpC+pafil/1bRZkgvKrFz1gM6TiO2p5BFJeLAdaRBto5XMAALyl/Urk9ot
ZlWaGsBo86PERScTy7wiiup9I3RJo687wvZLK90vDq5P4NVGXUgZ0YfoPH4EstwXHdxAfZTWubLh
n2SsLoPIpfKElXyBLrNRi/mKZs41PQSRmpsLK0GubeRcAh2UGU54+bzosMCvtyusmf9KhwyUmvl+
pQZCSyfPii4jVbEuW5w/g94+m0gda94y6p9eGW58xKWZrW5UmBtRyaiv4UeB192CxGwAVdyR/1w8
Y/C5ZKO3lPNdw4SyiRVob0JxENPX+Pyt4ZRITZXFbZE4IpZo+oiQfpO/2GhkgSekPFjHWZpzKFai
1KGNvo5llUJGIbdZ9/dUNT+67Ys8DhvpJP0gaGcPuYniU+MwajGxtAMxtOqEtMH/VUUEjtvXryRM
tzpNgkRyn3+oD7ZbVMV2pDlrRPOk0XY005vCkPiYICOD/x4j5LJjceVPySKExrRskkqD9AWb0kb6
hI22TO5hRbVE7DnQK/pIS4BtS57vk3wYa9+Ha/ir5TcdiCvlehpc3ioHWGcXLYLq0qnFo9ii922F
fTQ/HLstLN/c4uTK7OrNPmPpEW5Jsk6uIMa/22Q8QpdDBrXuDlSa8MEd7e6LjHypPZsR49fc3hZB
QR9Gn80A0awf0yADhabjJ+w00OzTcgqPJ3NWXVsdnkrhMV408nyVTLKvygpOEtgvWoegYwmTj0mX
h7GslC0zcfblc/RVQcrW9YDSyXu1qY1DSEaNr5jDxF0FoZOvxFq7qRNTaOOzahqwNm+tV4Ak24iJ
3jMzm5XyJ4hBXfT7aF1W0A6+5gDBH8sWyWxXKFQ8P5j64aPGcRYMPU2mxBbxMlkHFS3JXEaZrrG/
0cFrdnMwd6u0eEQSkf/tYDBhI6RUShpptOd6grs3TwYW/V+jvRraRKfQifpBGRKx1VkwpO4MkxjJ
U4oxqONei4HAJY17vyql1EtNidlQzLEcvP+dCXj3LyMISVJn8GD4tGRoIb9LBpF7uOPXe5m0PXjl
kNc+dvvfCEsto/bCNHsjIL7kRtOawMFQo5mAtohYmEGIzNum7kK2WjEApRNwJYYDd7OkxxMrQOIU
S7V74gJVI2CP0HIAD1UVmyE+aA14sVzSKaTxfHN7Q58h0KXVJIcqIScQQfG+vEZqOpQk5p83DmHn
Giw2yhNqDeac0x4zRaoVsSlMIY2E2zbpOwDHg9D1S1jkjmF3J4vAyZcHNjxRmmyycoO8t6lGh3xz
sM+007Q2t8PxWEETEjmlLJhtR39g857keOEQNdyrEfLn8CXvHlKiQlmbUaGk/9DURm3SyMIwBoxl
HyeA5qxMODewaiOImOUoE9O4WNxM6K2+xnI7qJ2TLHIRigDUVsW1Ae+27djL8GBcRWonaQjO9VsZ
5p7VXaC5gjg/DIvZrvHTv2OXUb7K+QI1w7O9Yn+iugkbe+bPsgcJYZGSsi8eNpnwnbaTAORm6dUl
9dqlFFtgbzk4uBruB9N10rfjktsNg6/XitekXzEtEqNTAgbikh4p4vEhj4z9jLpSh5nBBW8kfmi1
qrvfXJsA3NrYgJ4AygbFVYLVF/1SugYh6XdY0O2/YX+EKCnla9xaN2zfsWRcUzYoYd2fYZ4XfWn6
ijurZExRaFQi6psCvPFlif78miCeq2sxpSrNN+yVgJroLw5E9vQxMWFNkLnTorrj0vWpHZGaXeMC
DeYRdh/2rKf96bfOl1AW3cb/jUUUkoLVm7p1qEn6m2npNzPbnLV8oHDv/Y2OvkFpK7CRhRo23p5K
dzLFXQLp44uoI65OjyrUc/TuYzWkG7rs+JVPKfPNdg16xCwJNk80VolwQfi8sGARkvfqBEijoQZI
SzFBA1GK+6h8STJ6ugJjnhIoupsFTtF/JCteuYUYDPXqWJPmBTW6cKd2MPHTo2ZpO7SHZ+AAD2k+
ZUI77s0KxcQvbGt+KqhX7ceUE4c7n71QEWEiHTKhF7FT2UzdsupwkyzX3nOxj3FZJ6jpR6SrRO1S
prvT2tgTb/XkPc6CWl93EEh6xb+A2UEWOE1WnN0NY1eBVtRFEUqkUlgiP4NQdJ3EDsvS+jF7dI7m
VE26Ku6+FpTqtdOPATxJK5FvIkaXSYObR/xVAw64PkvCUsgYu19idkkONM0duWZG5vDwSWfYlNWf
1cTESnkeqz/xzc12lMT/Vw8I9xXyvsIrdbYWd0ruWO+c/aR4nmlBC6+AXZ6nskkhFASKI0QKT4S6
YQ4iVYjzdWZ9xP9MvX+PnGEhsiWlJ+ft/pUJNfYRzHNCVCB98Kp0/lr9C9QmbP/FAgKbQUbSk7In
WMdrM2unjwVYCgZ+wH/Uo+zfvIVUQEuS6PLFepBBkuWDiCv6UDv1qWwrhuR0Glc7EDmfweEM4lEk
+F8pB9GLIPhGNovvHKEU2kyw9Jj+r5ktOrtQTcNNNS8AMxNaARkh3psfysQhw4gz0vXejyDQui07
RIUotYEwtyXx5d8eLJUG4ypaWe9t9RnQi9I254KAFhdPTEb48+6onrIXUqJKCYD58ukegue5RU5x
1igTIGs9aBsRrnHIYOleIWasCsGzFhy3Krvnt1i6yiCXLA/wZxShYfS0Uk4C7hu6GygI2kenjl/T
wNOxxSVSj+ivyEc1tDpvlQP1EYcZagta3cMhmm4hdn/DTZULZMpt7FgbvJxdm8mfNfXiy8TxdDd7
CFg/1usk51z7Cmwy+Hap1VmOPgdBKFpbAdmgBVhiQ0LpLakXGv+hHHuawEs4CVeM0jIVyo3PmVYk
h9JQmVygb6NvBUQrgyhjv5FA4JFQq8iX1vGsoA0gwl1kBQKSd6JILqFEBQ0tlY5ffu4kE4kWdtqh
9WRDtOqR4TyxVkx6yDvEXGl6SOQ9uS/55BLctvGt8hWghhO1CIDwMmNEYKEf/GXf5OrPRNF6cQbM
PYEwAZJ5RcejRQXMmnrZ11jzicrofk8Q2jBJq+yfaNohY2+7j3SFl2p9LIo+o4vgOfgFG4C/78s5
92dbMM53qCxHFiJqGyIWNBocnDiCydYXn62OL+DFk4wnmVKRewmg58JsC4Ch1E27oBXk490iza8a
cYBbzOg9kMy1ugHCbSmiIzaJcEZ15EZEY4LHAuaq2SqS6MFZQNZIpgOqs2AuuWg3LWp8LFm0I1Ga
QBEpnc2CS+mMrpO5aEuk39di4savpD974hBIF7H9EhjXxBUcItRO/TZ3AegC+9SuNIjN9+jnwT0c
k20rJd13qNJ1QOSu92iSowPQYTTpdmsmrhAK7spAKgGMih8HvoZpHQ/SHrNku9PSshfHIg/nMiQt
DP3ZdAjxZeIlqjEf7jE8nit3ajsovGBSuQ9jj5csf045EOB8wdGPDa5RSOMjEa4D3vugWmPnP4Yv
7z8AnKbFIuaodH3ezaQSaLunn8etN/CkNHnHoXvGc90cfe/IcrE4WVtJAi9RnJ1669AdG7T0uWTP
KdIkpXpYyQ0AQjAQQKZ/jh6n19iO/Pi00cBGQTezzkfFMrgkjA4Ck+YojPIwjRI1YZEoJsxV1IRb
VCW82aeq/k+XzI+1gQ6IbDyTLJoYUz16cYIp56iyPXWXcYnZ05fJYic5q7e9DmyC1/30O+6XHIHU
hHB6d+B4FGkdm2tuGhMj0zcNU/ekHt47IRq1ANWXXLugObNoru5HrtnlhC2DGQw10lDmGyrsyeiT
Kc2+OuLBhmsX3IeQ0HFOScJCEGC5Mm1CDeM3e/VGqnvWp9a01qIQMontG98Y4eRDpZ3IbW4AaxW5
TL6AkXu1kALEBUjlJUraL8za+/giEIpdNt7vJ2rPLI2ORide12kt6CHWz5nlCpp6+p/z9KJC8Zgn
DaE9dPZnc5KYggEoJNSLbeCKDHklqJeLjIwIvucTpOJOfrPT02T33woe7VDMd2C8+Po8sLg9u1v/
61TRP8AvfL9n8sK3p6GL0lo8PnsCpkcj3mVg06vVCsRZWI4Fvue9hfbgQYGeKsQK3oFKP6w3xk5O
VOR3CAo1IAZ59ZFcipa4HvIkOnI8DYHZkWRk5j3Fnax6z9l6vVOmSmvkCpmmZ6nMqF62wotgFfi8
p6GFjf8GlGISQGLsP6JuVOIQbIoohrN0d9fJ1jarybuNY3ZgBmF0MFx89sN5HSe/sdnlDzBNKDlX
motc1JYc/M4pnlqDOksZ/6SFWY+k+reD/PBxkKtJIa5BfCN+EO47ZdGzf2Cfs0jTAuAm5svagxN7
2jqwpyZZkodEthSKld6Z29DYcTydfF9eWmpxOq6pPWStTk5h6eRTeKXKEarGWlvRUsixRmGsBKTw
GTmFcQc6R3/iJ0/BCo2ktRgCnI63s6rEXfz01HAsbW4DhLIs6dfjerTL3iSKB/1fTfB+RM6sUNUH
mW3xJeOXeArg4/HdNDORHknfnvPDKV4Dz5dMdm1r59jvzr3db7cV0rfHsPa3bNusTuACe29AbTum
CvymLnkkDZzCaFUR1oTnWPpevfuyYsyoDnXs9yndSdKoASAWjQdeYazn//00D38YU7v2HmueQgks
ZJ5P6PiU4VzpihRcNsnjSU8PE8ECGnRWudXOynjejXwkDjSHQnpVWUS2lQGm+NJdGKEOcnqeYf2K
qgRkvp+vVh13lJ3eo6p3G4UyewFd+2rgvX1IsLBJL0bC+gB4O62plwPFfesQ/JYNzRL9oPli0iiJ
GoMd5FmBFbQpdCo5y7nqIpBhqD0Tu1E9s1ETqvdATAAYC16GNiiMH2QgiA39SACcfM3jIbCcl3Fl
An94+Tp08mjhsxcwyOW9wb021W0QdfPJv2ejv0n/Nz/zWOiMurCxnBHgqBIjG6hDkvhjIp/+BcDe
FIpiQ+DuYzsRVMjDLmGjFV3rslwhJNb7bwAkDGoN8wFFjsL2l7FglimJnw6rzYJtmCy2bPYGC2Nf
xUZJ2BhkpK97DaIyJBp/Ds0c5Yr82rFtAg/g5CSHAn5tSdNudngjGrkD/LvKenbnnJIo5j1NFdMD
FkXrt2qS17ayknmJMPDNSo2VNOhUhOCvpsydQdvtAbjYeli53qGuExnbZzmRv/QdtJNOF1kxselb
m1yuKUWDASh7s4Z/TqpZG2WlDINssjDUkArfOC2kGLpjZbhEzFcUWUzZN/NtI7Uvc/pdMzuJEx1o
YMWRahNDc8Ve1MGEjRjBjZKP7sdEI4Rj3RA4Hmx6vS9XiIFp2SDSHYB0PN3UA5qbcXmK/FegxPXz
iXuvCK68xMJjNKH09LpeB961r4C74A8k188/2AG1JcKQN+XrmrxBXnCeFWaYUPKkO/JGcL+laxRZ
32Wn3kGKutSPokpMSttsYUAkucU5NtmwJusvJgmVEvXNxn614LpJ/h1g5VMXILpj3oyzYQcykS4+
RItaDkQysMcSC5NDi6jYkICPl2/+OCcujzyC9dL0QkOWDG08etyrKbmuGgjrbHpnczuJbafXrpMR
K8GImXgGKfPgm9PD60LkWnZde/Rg4vSgR4nZFLzCw79rpjBxDwLB0br6PRE/J3QfON7LtpnOXvdi
13xcmHnz6QUttq72QEmr4UAQccmepminj1qzOCQNHU7+WuhiBWaYpoMgtEl8Brf2Qsto8pxOX88J
ROJ+bwq1/sTm9qGqonyEzl7T+4PjDS+Hej3ug/eWjcx4rYlAS7Jg3lzg7upLZ7NnhW//q5pHY9PF
KsrYzTORBfd0GjFmrNG4yAG64JHJMIaE+VSkP4H2cGZDaLxgmuE2+6bbISrYfoCSmEkOt4dwfRqg
QDsSbOsYh36nHK87ve6oKJGKz7YPST7qeLd+HCvh0lBE9vp8h9QWgq1DDjlr73jji8msDcHtKL0p
XSOSsOXwxptJGF2jLy6EthB36Dqq2bGb7Yw0bVAOmy2RFqfe/OmVKnsE8JWAQaXb9Cj7O66Apjwk
nwxgvgXSqyfQXszBOb0HWEW51Ec85qSM3ioRUH9VBhXYu332gw9IixfMew74PAQz9YZ2JIqnxbgS
NL1kFFUI2Xj+QgukFgSvhIUsBouRK+8merFeOV/Wk8rJSIdrg8sPQcqSGxapKJAe4t1Irwk8gR5z
xJrahV8jAleoZrl2RBBKI3msP0TrNGa5+g/N757tGra4pxcIyAybTpMzKNep5NGa0rR2SiSJCwfR
9iUEEX/bkt0V2oJ4pLLyjwVdzvaA+EfulEKzo+NvO5SaJfGqpKtqHuPW423qyNCsfqu2Y83/OYgr
SUhvjvUycamx08aNgHxk8fPQYjnVdaEHsXdn7digkaqveJKqK71c29gbTIx/q6GclbIagluaCqGT
lasTN6Ozeke2iZhp2vKd2bzTEPrwRhPr7EYuXTq9DfeRFKXOnE3rrZoRJ2D79Xr10ExydtHghhFn
w65pySVM7Fh5klPc6kw8Ol4k1dAmmqJ6ydNFgoxLFCFahAkUIaPvR/vIzsfoKSTJyshWYmAhW11Y
L7a4odw06IKIAiYzToH5aczL31zTL33kvuJ8yOH6uZRSIEDo2pPF3pUTGsfj/YOd7HOAtpcKg/Wv
7K+LzY9bVSe+vgfgVnVWyADk3xeOyrmhPvM2Kz0BUWgYnowoVji7Fm/X3ssx3wXq7UpwvvREwjfV
0Vbk7KuYwntxuW2Zsdki3NjwRcGCHKBOMpg6UUak3uY6n4XrEb/t/VA4vI9UuH+crpCCx2LrIpyS
PNDvdaJ+DkCwkiQzSQDI9kMflYLB4ZoWdtJ8dXfg5hdhBAge+jRjX6sGUFX/s5f41saw7/Wzg9l2
qD1hob/W7MwPygxu+tNbpWkvylPVs1q9vXD0XvBfxhd75qIfFksRCGGKh8zTkA00J2/7ZgcT7LmR
7DqJ3A0OiMX0Q6g5lJb2ltVr7Qat6HuQfYxuXil68DPIh/HMKcIWr+LvhiiNB2ubnpRgXzJ5YhPT
0CiDbv/NIMLyhQX/xiPFpDqg5k6on4gXV+tVDFyfv1kYhwHr29/rcQsGMh0/QUE4/i+sSZOvaIrc
5WlFZcl+ZfTfwIP0l8UE6IvZxiodyjH9itTjjPgeZnzAA8VM8JQa+mLUYEZRUig2J34fkyPruT73
XSVkaD6pAPWNGv655EPobGjwrnEDdRHzfca4BU7mAxU/AQ99YXbu+GPmdJKOK3xNuc5oNe5NyXbX
lJgdK1f6P60lTVFZ6x2ZdF3ERmccL5CmmpjdUw23jZjj1fI3nUG9Zk+lL0HLMbhdt5FZ0PTEWa+I
ORrAntDVOnYiXtfbp+a3kLgm9VxCb6cB/xHCofGJmDi3AXIr8PZt6ls0eBuObpr0bLl/gHcXx/3s
1SHPsPu5mBrpOt7LBeX81nTvjjYtPY9nRt332pa25aUBDuPUF6oEnJw6UhnviFaVxgFArg/syaH9
YAnxFBiJvDMAoWdzmZzki283wqCH+8wkj8rR/6zttZXO/imxekchrH4Vd2KWMlsVa+zqlx6igN6k
K66szz/cEYmFbAkxmWx4Mr0dVy5waynINGDNi+rfPO6/eIEDw1aoynB12vRtxkraTcgK1t4b1Wr8
QQESoA4AXHxuAY1HvNpClKyiXZTxhjAqNyiEDnCXEliNlko6YmM9ot5eiAZdgrbmE2JjBLRjDaE8
XfOFFhoVT8Bylb7RPRRiX2fvqvGDLuXeEcRc33L4igWdGf1NMQmR4ZHPnv7rJXMNqDVAn/poUsUw
GyhzTESpIagpf+YgQ65OP/pFHAfiAZdn598ZdzvlLM4hjZK2dQXRrIQZWk1GNydqcjfOkPhYjkcg
PnYX++RhLE/kois5d9JbYAIwKht6KMWhBwVuzhzLeh+MFZ64KHQRWvigAtAcODP56/ccy0FjLohn
wcUJLUb88trK+76ILRJxSDBn4a+veQzX56pV+/Ce5OCuN2AtQ5/c35udesNFncUOGsV8/ibUtrBg
Ofb3BhiRYqWawr1eehhWvzwyWsubT7ILi2e+R49g9FFBvs9KLw2tT/5+jGzTKu3k5/CWhcAJqPQ1
fa4K/C/wcjqaxk7Q5uqW4A9CgpAj06aJzGouJPsWcLjctarGX6YOL0h1Au+tn0N7SreNQl97KtDf
yW9UhLaEZUanUG3978fvOopjagQGgALU1+X/1RLxny6RvCY4hgKSqQqvUeK6RGIq23NgJ4nbWdlo
r0HiPYGM0ZnR5R/PAbp7ZhUeouVwC6ALzAy98z07+KhnYTxDUJVbs0rsidpYFnSKgt1RKfEEE8Us
W2RMEeTKUw8fLqPP9neZYBIQQ4mLXezqTXAtzupgTGmasyt1G38w7g3f2S7Hu73nGMjf/gtumHEt
v39Kgpy4ZikBa2WwOPOV/J8wJ6WW5BbQRUpR6NbgytePLFhO/F2QmKRD1aTSzM5QR1NmwfKYva29
SoYiapxkv2B4t+BgmBle4ZlyPj5DenbYM8XzGvfFiYHDfGP4grlQuEM1ags06cidRsUFQCO+X8mM
z6r3mXgj08R9WwGDinlDe/mHezRXP1Hdvf6hltm0b/sqUJHFCb29tyelh5zdpwDKHf+DiO3iMqAd
51On/sp+fL+hg5WUO55md4s2KeLgB/EqdbUPplx1dfm5P069lq8VjFztztN3lDHvVPPrbM7lpjc/
oZR7THdSz3LY4fbKf42ccxFbEgiq9MyiT3uaPm5RTqrGO4X7oLyoNo/GkFuaLYacX2gddJKEOAiY
Ixx93B7JAwVzA3d8cO/cIGOidIwS8ag8fNyD5meZ8F3WdglI1gAoBAtzn9sbNCZm1UK8uKabgGr/
wDnVVN5mYyrbAhgdMc/AZd4Hub6G5qnivVriK4ajxEuWeJ8bykVy/qeiduVZG4FKFqy91FoTMZgc
5IgvTuk/e73/AK9VrFHjWWxDQUxU9K2wl/bFSYYnynVXngS+64WbTHEF3X6aiyBSmkO8vI9DS0Vu
YnSWDyciRaxN/iJ55ruOKgOIpLMOyMC0eJGTkPbTnwdkHw5+/FrcLaIVxWwC02I+KDjATswurhX4
dYOD8DoqNwVaVGkt/QhPP3xiK4SiHZbfrX46oYA75Ar7ut+nfwHVc0xsYc756vkwKSLxTZzjr6w7
TE4CrTTsnzQut2IFc8E8Xigc7Pa00IblZzGDFNNzkFHPjrFmZMaZzzMHPlfKzYHdarXHfORo5szJ
vPeTCnYmANt38v1BlWIrFA0LTyhhPjOdu/D1GOiPGPMXDjd3GCOCHWZszGfNJrQQwSkIjZ5tH0M/
MQaUBsbyjdFXPr6r8IE88zCSg16lLBdq1ucyCNBifbXTu9eEV9z2/y/8la0+7OCaih0hItdlP8+x
9+unCGbU95CNCyPjq4kHAPt146RHXKMd81oJdmD0CyiMjjESKZ1NMewgBOuDVk4Azkz6ECJfqQQv
GC88THBDeaQwv9F31HsNS4rWPhbaFxx8cHEKjuW21skxgAg1W9KG8LmazY4QGOLThChhMpZkkeOW
9cKeeC8VpHezep9oqhOfkALrl/4skl7zj9sjyOfNpSnoQQ8zu5UP7ZFh6FpPKT/fjAO84FhQSWsR
t6DRU+pfxDMPHZTsUQ8vrQ1/micXw9peRYXrW4ocfi4RHgdi/WB+yMBlic0fO4JGWlq9h1GVnAFM
4clHd84gW08qjqxv6jsS4ZsjrJUQDsSHtanbr5mKytizSjylm7QPPyFrf9GMz4BI1c4ShbeDS3xJ
1Yc8Wybz+POsJHET2JSqBbkOPP2JuCQgUSYxb84tQebEVCChI7XPNjQn9iQ1y72oZxa9df9SHZPh
yWWxfK9HvzvTh5rE4QzIiMG2f3Tp7T37p4dI2Y72l3MQzZchIKG8RmNR7BingfdA/O1kwUwFxrvL
kH+Wp58YHKDFq2CAA+nsTzG/4WE1Zso8rr/PbQcy2090EvoRGFUshI9biXT95i04BWhzPwveDv3B
rGs05SlchqwebMCenqX9ZT+zKc+XKdyIVPjzmCfRvPTmAzogIGJ1VdOmVp/1T7vPSxV++a4Ex9kQ
5YhNl3zhcIbya30mmxctqmlmJ6QvNrhi0+x3x8oCk9mQUpEcksgSmtzYd4Wl5NxhuP1RV66sSGHT
PQLK9HzsyUh0GR456LuTN7QTQx5NyRyfS3CC1+paNa/goDC3/tbve8g6xr7Ie8WE6uRoiWFvJO0J
5UnSFGQ3G7CYdAM1YIV5oUX2J5LwaHzg0iZAB9V1rTwJxTG0mAUeVM4CPhQEWz77f9Qq4nL9uP/7
YZGHbQQ3VsG+mgmJ+zP0TAXGcKKuCvkm44vbXwil02nck+VFXKttTN0hmGYwXxoIQzXd2K4jkMJ8
3XGEbqwQdF3D1l5aOKI5tkTTExi0fqCmguj9wIRSdenJmRQKrrqw/0rkoSmTw2tnLuAyWG+WKzir
0O59OBjqyKe6UkjYgB89i/Pyec+ead7h/sEZ7x+Zki9YByMCSpB7rgj4dDSKsO5jYqWA66RWv3Kw
1i/xY1izxuoB0yxOf0aQ2WkRXMmw/XaP+bJB9svwbuoc92JPdkZDtbihvupH0g8gq1m+aNoBhOv+
CGJLlBi3ZCaUHb1xXeRMi4sKiOzYNXqaz0fP/I4msbEWI/8hhw6koL8hspRjzj87ie1UApr0oaVF
Dlvnb1BgszjR5cw4WVkndfSiBuD/N8izd7DhwxyG7GyozPStBljfOo6YB8qhQavzMVr5mG2bYfik
BG1JfxMbwM+0xjlo0cyBAMfqBawDua6x8j1uR4ecKPzudckjV2VlZ5mkDjLgNcCyR2BMO21S1Fd9
1pdASZYNdSfZr8PTRHitAULsyvZiYkIutiMMJOHY6qDThtxy8OG7e/hioGNG0jFYgumjGnNG6iU3
tKeB+vqxlKNRusDIAWTeR5zew7BpsP5zE+SDPjfRd1vGnMSmdM5wT5GXvp0cPJwvMaQ92kulHq7U
/6msRO3Puc9CPpZo+4iAy6KVqF2QBaN6hQfpeG7tCMY4Fke0kxr0GDHblDBkRoXOz5FL1hmAGfX3
8F/MEQkXyJdLLKAJUvP1q2VOKwVFZMM5ObhEC3/H9DxxaMYDthQEteMYMHUALK61ABP0YfVtgZ06
lnTXxCzI0/Ox1D1g/vEexqV3Qz7xJCddcBrGC6EVhfvmeBVa6iPRXwHueNPv11QuSzSDOYWxSwTa
jSTjNQGHjDv1MrPVoU9h2Og9iA+G5DG6zjdqNa9cdciwcOFUCYgDdBrBaXM2cl3TZGHdAyid+GN6
6jHsSS2ZWSgRhmfatXGWteGQZjZolnVVgdfdbqCmEiBvXN7LpZUvSRgurqX5BmAF3OA3xbfs9pnn
gt/N5KMk/Vu50y/RRkw2DGzJmmYXpEdyBVOy2buxKWd7hNAlMl0fY2szv60Ws1Vy0awTZyOZpD4b
nVwYIH5Q06/N/tZdQydFfy6jZfcs5GqdBxI9cg/SvIwnCurB3PHpWF6DH2FF4hVg+MsqMN/zwg9D
NfwGNuPboIv4w2CPbK4zGdRDwnfhThwP2hc56o6IDv7hwFDmFZXOSzyi/LBnKzvLiFEmw0GgRolM
ePM2iXGjS1t1wDWxm74TLyuSPc9uqDS+/oz7H7SsGxZA3AQqC017LyeNRzBDcQZr7t40nIH/ovey
AxJsLF0dDYqJIvi1A+SQso9iRffmo5l44pp4xDg/QhNHmE8gmVHtZpeSjqgjPgjtrrnGwA1uuYao
JwFgYJMMx1vXb8XXi4EY4bsVZxK4VozK9r0v2RZ2426yqas4rZ5/cju83lEfOYTck9L8oj75ZfBi
Lhz4ljSISN5k9MiQ+KdgmHpD3XLCaj0IY34G3JOG3LUkNIi0bA1furzl4fInwAAf5c88pTzumpG0
mMUWwjO34Ntd58O03qrIIDjm0jOYGAsrnMRYKn1SOOvNtDzIt+2RROJYFNvvflkAN26p6hqGoi6g
1lijmsyWnCzL15AaqqMvZze08lT+Ctm65o0RvMGlCeA6EU8Xavy6nC5vEf7epPDbLyKCHgcD64Uh
5W/VvxdZa4hPJgSmT4mCNUEUe8Yj6bd1no7b68tJmgJhDig6hsGJl610DgbcaZNKCqndUjcc/nDf
a7wmDxUixx2iyChSt2mdTz37ViyfuF/04WzhisaXqoXsxQQuTFAMtBepIlkIueFON2+AwWCJq2Y0
WkMn8QN7ZILK5NW1VHlVxCwSX7jJBCvdn9XiPwFQYlSLxFy4m1jjdhkogLJbooD6aQRDFauX3NuW
YdfHqZ4iMD7t/dEovM0OHp9efj69HP1WCTnTTnCkCzaT7KxKvxgQJO7mSgyjaKQuELc9E9D6krcZ
WOmkpUgeMeVzg/UPnlsE1Tjk9A5DyXOX17tvYKknTvRNCgtG+1XPFi0q9nD+63jqgwuHUZmTTe7U
60V9u/m+aliq1n8ojq+PSMbSMuX8CCBbw2OrnWCmDP32qS6ss6CK/I0gED7sw7TmRWsYoYhFDH/U
jgG4iIciSQmNkhdKN5iGBlLr2sB5dRQYe7c3bMOLlDGYV3bqX/YQPs06ZVLafATRt1itolZh6NDo
zs7tRT0vlEmO7E3+Xm+EzBMtXtfPQGGSLpBsYyMyt+BYOxeVeRmDQNnqcaLMNY5jE2q0cugmqnUE
X4IhTJJlq+RznhLtnoESPwRF7vbcDvluJLuaYlc/3pdLiVQPiU3FRVXaYrQ9qWMeX0DieJVj+O4/
/hK1iviex3FxpZUAmlTzUP/ELQw36MHcVluqVCdxgNCkT+Bg1Veh+tfCguxuZHje0Yt+tmnftZPy
PT+hHEPEX4eHxeXUyuAYiDnnc0tC0NqCQ9c3HZ8Fqq+QSAWqM88SLeUILH5hCLY1gE/vAunENxTX
sBYhz6Ake4lvfQA+YEqfAkxfugNezeow6h4kkzt9RF585jo1OBVCfez23yp1v+R7Qa4ZfXBZZdF3
Xs9+45HPgu/Xa+hKNkD1vSWHka9OxE+69IhYQ/Rs2/Ph4CHpOkQ2l5kkkCHbqXT/Veu0jz15OwBu
UgEVc2xyCP3tt91Sjm6AoAZ6/CV938Wvi89bHhp1B9/AvAoq/MZrohSMJ5oRj3yXoWXicVLOb14P
GXC9qvcYaHfzl1U+vVvUybHeWrsbPCGV2t0oaFIbMZkHsbWQZ8RCW3FVoBPB+tF42hdszkp8zbaG
+mUNTlLnRdVQtfXeN5E8ESYWITXlUUrornesNaZhCir8Lm9SuWBsvQgM/ZXPMMSx6y9t/iOdlP6c
BEXQ7JawJcA7KBjav3P3GbvH0Zlp9/ci7fQGw13vDmqnSQ+7Bhg2r+Y3SYpIPvPsnEHcmphv1Cgr
EZlKUm1P9tWcQXTjcoEB71aVTfOGeZTbbFVcrNgFvHXpRFL/C47x7VPRq95wGarezNCyB4nytRAc
+fZ/1JoJhqfOyQIWJeNfkK+eGSYlNPHMbQFWhN+o0/4W+CoubTyps1IDJbTvT6nIUxE1utq0d3fo
W3uiUS1C0nH7SSFemESvluzvrefu+I2iGRd0pGheAQW3C3VXNMawYgk+IdJ3GkC8gj02GYQ+aE5a
AwvUDGLFxa/L5w+nxtQpLiNQG3TiuNgRt4zq5JudzARjNRLwfWekJ/91Uo7Ir8mlfrFoFrFh5fFE
R8I4DwoNEJ3ywEx/5wRo2/g8MHsYUpPfp8Ky2KmUpLiDJN6doBGbFIhXGpMisVpiJSnitrk1bPFb
svAVsHrXD6aH1TPntIZngJM0kTZ7HpRwgWTelBuEUUu7wc8004K5yCA8swmph0ayBNRnC8FDDijD
gOJnFIKA6zFK+EtbcPDBQ1mVhAJbpCkux0ld667Y2Go9tYFXiK+WWJRO5EV+kJyPrqxdD2rhq7mj
RHjdea34AmUqXpRLZVOTOl9CbMIL0wNvU8Z83GHL6cXscgEepb8ycwsMRHgYJApIHr8/f1cNRGyf
/Fm5M6P9FdSTXAUNJPdKrni77d8nsvpRTwpF5I4Gu0nxW1YS2U9YjGjk4zbnR4wJp19oC+TTXHEB
khZhcFcTOyD8mAp+N+B4wOhp2+W3rSMjeeDV2c00Q7Vc71ms0RxmvoFgb2yPMiTJ/rFKbwOQkru6
bzHb621PhB7fKEAiHrtfOcKSpBo+XhOLz+2LbJqu9i1vY86kZHOYxdMy+P15I+UJr0q3edHnBK8E
4xtgmBOhaW0i87nfo6mfX4/XnszCUM8xOiMBZH57qFHTPfa/HA0yBz9dbAB+dvZ2vQ1G2G5Zlc+1
sKIkyCTA8NousuOnpj2gBWNhmoXDARXo3w1YLJ3gCTo9T3zw0nM8Pn6NGy3M26Y/7tUPx/hTjaRg
O5V3cACUCgToeAqLPWT0Qgd/Tgjh9RtHklKQu5bJ2nZSbzymwK/ZMxUcMFJYAsum7Z/RL6bFMin8
BjozE6o0Ip43aSfuj0VUpLZo2otKzlvQww6Goh/zMe/RELakMTlRRYx638c+Xq7qrn9OWnrGLiCa
TmwG5YYgW/pDBkejkQcZcf1gh6epEoKQcwuWljs6BT0K8dHBsKfiS4EZ3pkL62D7WtNVhrT8uyj8
YgttU4J3j1oU12tJoxEi5nakrduK5iqk7R3iJwZLhAGfhSNLYzPRJVApw/pvL4EjFOWh4p9/GCzO
C7Jh8K/2YyxOI9Q0k9FMGDjgcEYG6mARDmgNBqraGSa3yGjxirgMjMqV5URzQDnkSM80qx4NHDLR
ResV4pbbrAtaCWb7yD5xM5XJsGf9opfKOF7nwpuHQMYG8AX63n3DitqWSWB9BE+AsSj/T7g2eDqS
9cMkAnGF3v9OOc9GRue2jG0d2aR3OvBI7zsRNfZ+gTycA3NVJN58Awmh7V1inMplBQ7279Hraz7b
BV+ahsEhvmlHfospZwJSQdi9q43TYrVrVsKkd5RmYmjV8ABDqCSm/XUSA/X/e960yqcBO7bAqFSH
hO/37l/xkMb7CZhXn/3/oEu0IeqW5KlCir9w8IuiveB7biYx4gAp7YwN2+ttFxPBWsa5EsDLTNQO
VjB3onwZN9BIv0DY0FPGA+CVf4Syn8M9yrR/rNYypXg5n2mZkKgtbIFxWtrG987vKIb3aXdHkq2R
X43B1UtKYzoJPKQAczsS+C82WgQHj9eye+6Upq1v20npBGTpBYCOIJ9Xsw/y+w8EtTBKkH1up1ka
9AWq2i+waGVix/lgrQYOeMKazde7QU4E/duMkYCVvAFCldrcb0m4nu05HI/2Dq6immXQY2deUV/h
JuZqOzB0lzmDdY8rugkpfxLN49Vpe4GwQjwaWezh/6CMlpp8Dc5zV/+0dGNKW1yYQEKDZGxwz/ry
ZeF1BRefE3VLQXZIggjDsymD5m/veJoGA3yk7xeh5gBwIdpku/vtneQJT7/IDkYrtlfrQ2A+lvt3
jyMC+tREOH3u1TktrAOA8dS+skhhcq0DOVUnOEfKb6WabBE9HWP2OVqRG++MgK1sHUQ4V0TAbb0c
PRLR5+TGB5FapH2sdDlEFm7jNkGOVSsBokD+Yl973hfLE7YMEA9BJtCKEuhPxVOwazOHSbjyCmKg
jMk36zXCKrNqSFM8coSFix5j3ehHDiWH/lrxowv4GHARv8cyQCFscmEHEozB+JeFvA7THpk+reyP
4pJ7COjt/Mex7gI4Yr+kDEqRg1ErLUyU+0gVPEbrxUL4P6ELlpIdFZ+7+sg5eU2CR08cMaarfkFu
mzPBLeKNor/uoeuSYPv08D+LhDoR2xaPWK/i5Ff81kL57XoqE8t04IIAiK/UdQsnVLsJ1NiNrrHW
qrEZpcqvjzMou6TABSvbkFYjH/zXiYfHYivZGmW50Uh5LnodgoXOu3aWNtGFkHcGBk1OS2QCoVtM
Vk9vQ9h422DIRMHLKkcns/BQqHoQbzNLYVWBSoFU1/bfarhvcQFNxEm2RibY2ffn8yIQlEUNR1AJ
CzCKdUKaiim6WN2prk0mbHhfUVS5YAMRiwIydczKqD+Xv5FEsYPupbkP6feDnWCev4eca4Z6bqG0
dpw4VKjTFm4k/UaywVg2r3V0z3J7D0S62G8tQdk0M20E9fF4stpfXrbnGsCsH1CjLIIp3k+ugjRC
x2bJ4v2xa+Ia/SxskJ25IXdMjaOzLG1bJGVw2P++o5b9uXaehINwlc3E7SmNUZXtcN1hAKUObomX
U5vEb8Euf42C/1DCBkw3/C8ysuXMioU8P8SPchjfvF9nxl6NjecHf9y3l7bN8ZXD9QIXlebArZj7
YYa5cBpmLze+NG6b6Ru+PbqbYapI09Cj15teJ2eQc5pCt2I3X3VNBRO6I9oL2fzn2rziwqKiLAe/
w09D1sOuyWBi33A3ykLfcDlxjz7hyvaCWn0RCM92+d7fQjrBIgkVRt/O2cO8Yi3+yy0gsmGNKJFi
Gfd6OSCiVLdqNYRNSw+TgTiduycdbdivheNDDS6q4dX501yAr1tpak6WcmNEr/cv5Ly/wnpdycNr
dUSKAtOHA21YIp9Vx7akgUaELfvekm1qOeDvTxDLgOyYeXomVnUCIQ2HqhkUUNYr6TsGOJSrEpFc
4lxeFMS42jczVWw7ZPt/yWsE3uvc35CHfICj/L+Uz5PkPuoSIddDz+9N3dE4Xp4rEF1UTCKMODxw
RsOnOxTCnpb3QDwCIzFy5PRJQG6ZeZ8MmdX7OUb1eEmAmD+ASMWzBlk76JW4Pzh/B9n0anHTYolr
MCgN2ZFfJkmKwZkO7DKMGB37dRz6WZQNFRQViMqM56NOkBXpwbt00nS2mtYqdzWDJDThAAuRBFMR
WENqtn9P8F3vX8/VAyCkQ4BBxFzr32o47ZsKb7Cu17XDV5VQeLAvZcZCr6/vHRx68Pck0g9o17xq
mV34YIHTU9ij4NLjNhl8l8AkaO0lN44M5PUE8GgYnp5pfstep1RmiVBznof/EgEkiC1Gv7GAp4A2
wG+kEygvNlBj3RAEGfGzP8PWkP0X8Ue62C7KfqS5V6IrrLZ+xaeLL93i7DzyjOleyK75qjB3yS5a
QNabGegiWYBvLxSDoLAbt2YZkv3eyWKIG7nyDMMqNTQpuu43v3RUlcuoCeWHu7sUfbHimQmHKtJ8
xBJOnjCs96lUHSTzG3Wqait6PSxwQVIeXha78+y9Fn1Aoo6jkEkZLoeCP2QHw24ev90kPGTgWZnA
1yxPXMEnis7VoOf1ALihy3Dli0ilg59lh9oIZ5G8wXMH8Rb881iZzJWmgx9AjyQO52Pr75Nq5r4R
UF3ImqdmRA9OcYPct0p0nNxA2ZCnMEMOT/2fno7qoKGDIGzXgCllc5tDyfAqJLAE4hX7Jsg7Grw7
jP8mlD3Hz0MyKLDshDRLtjxxfKBclQeLRUkJaTOdB6hpebBpiVW6U16eRty+nXZeFdzGdj4H+LVI
mV+EG9A4dbqJbl1xlD4+u1YBexJHCtEvl6HbGsVqwfA0hHkbsiQeOt1S5n4CSaARvPmy/cbShcLT
4Dwsmf+J9Jb0hu6EXIkh/hwil9glC/3nSx/laqVoAD8s080llZlar4oSTo8syE1S5DT6g8Q7r5Ub
MXpM4exXPkmL/YH/gUOGEDfUsstxaR/vtwd0yPtGOa0lMQUFEhCwjaCSjW1CXKMTc9JL1K4caMwE
Pxs5qSB1livyi1UoKifttgRLq/sHMBgtZTsGjSNqef81CvG0G4ebIh7bPE8FsHWR5y6i+XbGwULi
N/umv1b3Rr5Y5EsQjvquWegg+dHMaQxKxG6S8kt7B6EDokyoAxi5BluE3Vz5ERKAfSjlsSWbDOcX
WazAlau9KH5qg9tWljXcTZN/D5C/uh0FYtXk2H6Z6cgPY2rSpj0gr3v5KOW20PJWYxhMPt3pY0qs
UWD5eknf1DaKOlq5eABAeiUACB2c7rE5odbJLMydSZhtI0Aaaj0vMNubYM2qkGTHgM8VlgbzDIQ0
emw3dVPEitzLY5UdRaoJmEnSDdtiZT8wMTYwdiB9Twg+8YmTPM99jEg4yG9SpDGG/U4MncHpiByt
8ubt6+D36e+N9BuGaGI8oa4LUc73S05nNwuzjD4Fw75br7Ag072N7VThrlTKto+w7UEInBxkKDcn
QS1VtR8hcNOISMBkOyCUZu/XUIqO6zI/w9RX+f1p3sz89z6xjs1Hrt87juzpANqHv7GPbuqCKLV/
o792K4kQQyPK+mA0JhwVQvlgwvytqRVx6YSINrLW/k+OGWItqmtvZWsu2B9ukVUb1q/cAHWpHpBa
QEEwa+ePi0hrYgcBYo//BJiWkT4PSLi4XIxeH81WkCyBc5LwLU7vVUbF7fFFNgiED3PHupqawb6/
M+Y9SmcEvXRXCNDh+xHf7lx3Y9WWGDbAVxq0L/E382gvCMrJHCdcVjwz9MzyX352eXJL1aV6vUD0
5ogY9csWGqZOgcUhC2+QlKbuQ3H7QIVtBVassmJKlj03aQGioYkC8fcD8EY8zUeeFl/akgrVZ18Q
mpAd4VQAoulM6r7DjqbqeSrAu6+3EcxRBrRvXAMUL9ONdZa858TRN9MZ6XPMziZF35+/mx/jY+to
SpzDU4CkYUvyHOH5FJSaJBSeo9rf20UrWOUz/xJhy/KoMOWh+rFCEL/G1CaBJkVL4TClgNifOuJ3
ILF1h4y4hiQLEC/tb5qVBDt9kCacXZ0EGjUu2AX1jPaA9zvQWA/vTljNxf3Ce/Yv1tEoE9/1bX3k
0inuB7opaLfctMFV3WSMPnI2y6hEH6FlkdNsiIoib+K4U9p/UjANstqUV0huT5qQyZ9zob6YY4OG
ZccCfrXjEDA67hS0ukvhnpfMDxkDzlJXZXkzZB1VJvy72t5Yc5k1LKUw0Ioih5R+vgibuvaQNVZR
olj884DA0V1rHSoxK+DJ95T5bRcg/knhLaVR72hA+WOrppIiqExrbgwKrhzyo3cO1HeKtiPbfXhk
BbcE4DWNm8kXnpPdhvOl4/sZC4cYeta0GGDgwH2m2H9/MmIFGEIY18r1igOxwmxRMz34Nve4/f9V
YEmJe5mxI1SMvfRvFqfdKIbUkbqg7EaKiEgLdLQ916G5HyyLZhVsup8cU6HLM6pF2jadtHgL7V4E
m9R+wIq0LWTP1Cm7v4keBGBf4ufxhBV69FWDjHVYnyOV9W8jKG8CqxhNRxo1o0Nut7efMc4AesF1
4npzmMJIeYaxhuIgoozerbpNEvGTBYeQzeICmPzvckf4e/m1XLWZdrCa79AFcFqXW7ZWQ8sXcNyI
9YpXC/6hXybuC8QBYGQcHaASfJ/5JcGBAluqUArGxm5wosRC86S5Q87BtUUF4iF6wB//ifkHoftH
WnsB8scfHdCjpGLw4MAC4P/iSJub2QTtZoLStTwmuKOGk8/1KZeO5Dy37nlKZxhNEVbXWvGgEwVS
SqQbbagXx5lrVK08vMP54lhjjv4ntBhxN5j0DJLI+iAtB4GM3lXyCnuktI/GWroppWKrQFBVdGr3
0ZH+5kI5OdeNE09bH4RByeIA1Ehr4l0Lvr66FGNR8l4fw2WdU4phG89VvzRerpAlu6hjxLH+3/ur
lyeLVURYb0JitSfv7uBi653jmJpDR7ePGZTNze7ocQ4MDWr1CIkSdBuEcayBU9KwuJ7y8KyGmKbt
4j7DrVOvUUO99uQL0QaaStJ/ZAWj8YA4bFQYdOYcMYlF4FhrdwFMer4TmEFcRPt2jjDFoHJPgUhd
Ioe8y/8UmlTtdGli5+8/YEQo8E6uEo58wI3uCr14Bf1jqdzM3OL6d4zP3SoXBKH/Wfplm0NYHD8M
i2Zmaa6JF+DjkBvzd0QzglkksT1qn4qVI7YMUyX9QGRl6yv4l3VdEHM+R4z1BDqpdRY7i27YjqEf
PpYp4k9lZNoAcqeuy0IdOe0Ep5YKYNf0tTy5NVpfhBHF5cPYcBMyWddVSETqrxR7myeOTRE6E9yR
gxWtuZFqltUObQGrlX2PMwJjX5OACSVGh/QBeP45I/V0DCURwproqYUl7bFSjnsfUeAfX2GT09x7
S3DpIjJRasqJIN10/y+nkgodAI7XBKL0JvhaEBb8Rb1FUyw0yVzWUccQO1BQJJLKsAJsmj+5yEFo
hiDG4LGtNnEFkZ3vc2bmtNfUEwYxBlEnhqRBE0TOekCQOlS/vBqARnmtr9y95fi2zHBi5dPvjeMz
0xc03P01weptaDvB9rqHgcbNH11A8GTQDSaI+YZL51YK2nTWu0hAS01E2Q536zi2/9nWYGpvCGP4
Ds8K9oARKf6OobDhJkWC7wN8clyEPl+4hA80LiHARvEn/VTfJiuntdCE9OLCDzR6A7ITtC51FLWy
d2sFNp06Fj2Wm/O+IrnpIoDBKeqDkbC+kZJvI69KY7GNU0T8tvSe4Vlq25zMCy+ZizSPFO8cvvgh
Y84dDd2Kfzut0E9lprzF7vrLeafCUN2mGyW9yNAXIusGmwXLBvYP4/mIaddP0DU0msv0T+65K+c5
bqwJ2y0aBf+yljX9RRxtf9FwIckKxGh3v9iQR7oMNYuzYheEzpniyEeFYU93cNJBqDmgLGgQYf6w
k5fpwWmw27BFlhURxl2S9maJwwVSnUXNrXHn17QiuZ/yTNG8pogOxmb9FNQHjjs4/5o1vTCx/8Eq
CP+jvPNucHItPaPYIJbaAYp4fw1RZmQrfntBwlMWn7tEictiXYNOa3N+d+P5h+TLWa0AM25K43LS
2TyZMPKK7WP3rU+SRHocT9di17jL/4H0uW/6Ygb93ImSYMIQS7iktuvlCKNDzMjXdphfImY2/ChL
eitbnhmwVk65bXHFd1VeE+7Ex3a3DPPQhxH3YTt7vBH7Ck+tqHpqJbRu/psAFxlSFkyCY0O8ak03
vV/PuVM8e1WXgL5f9J1xCRFSjNNCdq/+fc8TfLYVEjkK2/5ViHDfZaNOTAhgmn04kpbWYCXIfxdz
kKZblCR5gpQxXzI/iwJHeW128IxBQ4A9/81Kn/8n33Pvm9+m9Sb/z6GgSBUEBZf8FotDZUl8t/eg
yiPSIbtap5GfNqBD/dsq0OHXR6kdWsTg4IR+2aFqsOhq5YKRTvVdakCGqIaC1VNyUTuR+/ZwiVGr
JEJH2xjK/YVTB8NWigt6ERJyvHePkJbzfdy5lxj5Katl8Gte0pWLMruQDExmYJ2qtWw/2+Lor7SH
AlykeMjiTk/Mb0h0ZM3FRNBoVcfhPxImcnBwUNLVfXMatFjeFkt/fTS14ixiB7wKXn99VpEYhAGK
D9WmVDA28sWJx5jCQw0Eebe5u98UWnrv9i8EfXlxTcZuxpUPFqGZMoEd/pmjJ8BIT+HnxXkzr8xB
4MuygYaYfNruVJz8NeP4OP/oOEPSnIwlGVLqkfTvS89GpZlHuabhv66bHoAF2Oqsbrgku2bCOibt
ZZnY0av75mAGIM3Vs/PN0CcblKF+USuroouKAju4elVbYQE9ZLHdE0+bac3mBnPXnxXey4hX8y0k
hUS215I5OWy2QaFX1TyrrQqfzXE005dy5KQw0bZSBLIItfAH+H0n3DAEaOx9IX+eMaz0eJ0Oypfr
yKVRP/c+Oik8MLzl7qMYn+up+DAGMI3uNtdrmXnzV/AF6hQ+rHTiPOFS3HpuGs5ngJw0WqNbLLCE
JR7ilhq2Izg+mtFyxyhyVI9P9Mas3EwrMPvqz9aUE3vlySfzSawmb6psWBio2ujiff8kzXmKjmGT
F0lAzvG7SruHuw4eIX/CHZM7Dfgp1xq2YNthRblfO5gl06d9xCpFqY9Mw6QkWKeVuuIJXGcjMb7J
dNhDfMrUiAS8xI68QVMSWV5rS2Ynys7iPcQG7J+8kGJFyBF8MRZS8kYumLPzY+qCO1lbVUdqBdoK
BPH3oG4jZKi/uhnHQCVDDjOWMp35XEJJk2QsduN0P0nSGJSjM679tBdpLzmVpkxvuhFeXNF3Lx2G
mkoUqR1oTPuAWRMVw/Nn5JPnmqvk+sCvj8bqfOUT3q4jtRg+YnGlR/2Zlui8FW27XN3qRNCVGHPC
Nj/qsX/KpE7nRqhlSkDK6Me/by3zFqQhbiwanushF4tGJvrSzC6vJxfg4xTEdnWEhhBDepuJcoC6
Diz69lN07L8rWTrGD2PaAkcxUXFtSo/YgdKshuTZ0+u+nLHX//IXYB1meFmoSNldZrOB4UGK4ro0
sms/sL3sp/rCrAGLuPYLWb/p/6TRW6kTsGGWIBgvydqwJK4V6ysVj+465y1qkRi48/vhqe0Nle0c
/05AeNHU6Typol/88IwdPZuq7teP54HwWabjlL+VfKkXbPdPhkXjNrzExxbfCI45f63/IuoXpx5o
mrdO9u2cFLrG74efSG+9kKf0BeaQsdswZvRtT4YThaYai0nxaXPxED7qyQFwLjKjyhewWwgEVzNe
SdliYDRDkqpa+D7wV/Ryl+1GXMrsXGpvuDe/WvArJ0MSkdN1hlTzj4yuo2jHZ1PoCGGzWFLKrQbz
xVhRlyVIcH3jjvoeo2TM3s4lMJbftK1tJogDUl11KVPpitdb42u97OeqvD7yfQq096EYftC9BiJl
G/HY5RsAZogbkwnabSr9jpZv0tbjgGNk7NufZocZru87t0478dfvmfiZLJN5ERqiwcvY1O+ikdRW
5YlmCKmO3plsBnVjAtO+eZzvO+jpZ+m17gRh62F8a2jnvCipPtTIDxYwvhLyZGmCzZ0FtycWXMsC
6eo6or3EaJrlyX0h5LyY78Yj/PWvAefGAKYGp/Pp7LxhR34gDMNekvWAG67nFG/iHvzVvFLoIC6b
gUhawXRRiPH4KqXAUmplwChTc/cZ1K/gc/j5qxTATn/W25T365xq46l/kqOQBXj/h5+463/4g+qc
PhDkUlmMPWKw1r00BWt2jrG/c2P0w6beGi71jXzOpdQdlbFNV30cVh8HHu+2JumDAl9aUFVbVVK2
E6j/bjJxFgpZcomgPmd3UiS325qblK2aOCe83CaAzcraSzGM0kfX+A9VCtz8Dv4mCGBWgU7/Mc/V
gDXFtwiPLqJfj8pEWrAgxwD7fnHhEiw3Jx7JtdFmOYUJzWbmOORH8UdmwCy+EHbDyCYKp3GCPfjN
2M4SGETihhfVmQ8Xz2oolUIf9b2H86hA5xiGhpb8wyfRUl4OVNcFHPJOM19i50sGXqlqjUzjmLg0
DW1IvH/6+v0aSE7NJMyuz7N1s44l8wjgBepro94eBupYGSnJs9O3tW/x/B0cWu901Qthxh/Iak8W
QsR0NsAsWVyTSJuEiLoiAc7i6kPvQ66ArSZN+e2t72OsIR2fCFJ/fJgtUiPHvMVpMxSCBdlFCRWW
wb6BtwLl0NISPS32dHXE+c8KNkoyXo4Ko1S9x+/fPKt2w68ML8SbvQLhObbW9yrUjYZjoWgeJAzF
hawZTbDDrnGKhPbgALb81Ibo3xsXWLdAx2p+fM3pBS2pt9Q/plBLIa8/tBPCno0IMXSpH+iSXUvJ
i6cvbJ/hvqIC6hhWSAbHhL58l0SyUae2riZRLhU6NwgdMJTusOQxX4PL7zp/0UVhng/3Aqc1cJjX
j9cHGCcbUUfbNyQpUpUcDV0kpCcoFHGWqCdXf7KsQyCqqbQC7IGx1Dz6fsyifCCHrPxaZpCIclwm
9dSELJ8sVQJWGg0329xR5Vzo7k9aqQn1KKbqmOluhg/t0mbbwunTw8SvuQikHZo+tcI3hkLRsZAI
jvVqdUhiAGEKYQsDSc5aygCbCiNwD/24VAJ3FW2MIMZzdqZAqD3972+Ry3/zqM5sC5cUOo+vmsSv
JA6YxKkYRssR2iqlTxR1mR/1LHFaYqcMou7qyWeuGs9QpeLIHl+ZUK/1urwaxyhs5E/5vcxm7Zfl
FpgAJU2gnUSHsWyqTsP/et6t0sfH+awC3mnEG46updHyUVX62Keptry6lq6LICLpplR+m7O1kzdq
khKyJFrIMCpUmNUaX4yofpjKxaNWg9Qj0494nJRyYelQqsSB5fedgJS0wA7O977TDqILk+u+ZX69
ijXzxTJLL2vA2zUafXNHEmahFbXAsRyQW18C+vUePYyyZK4uwPXOjwGaQj+GZAS1cD19sZwGIjmP
Kx8VoUFFhnsjrmTSCXT1NXaJkYrZsR0FKPzEI4/eLmusD4RCEz/jtwXyp9ZaG9vlg+Y8Z5ZAk3g3
S64A+w1eJ7+fOIUYm2AHxG3k3iCPAe4Q1CxqqOmv7BQQQ0YARgp27ZbO3FiktgJNJLRFCKygHP7f
5ziKWxA8RAeGXQN/VPgPmTWYA9kGps+Xe3+WHpKtamny4UTQqDWpapdRFi3uLf3tj1Lp2damMPgY
EijfT73fUxYRmMI1x8R7usSZaBwfhg/SNqMoTNlcgrDOOqfLw0R9E6Yqr26aPAGmvbGpz0OsF8v1
VWNeBzIf+FKOkCbI2gFRz75sTeC3cKclVUYO8EaWNUADaH+ffpqZDkJId2SMojrlwXVncVl12XsE
Aj0nZcmuEz93RoaL9w/gb91e3xaN0sh90ZGQkx5pMTuekdUy48O0gp8WK8iugT7f6735+lAc8CMB
mWGVS5DPZEMa74j2vQ0Ofa8AWpSVYo5Ey2MQMtw9BLJUboVErr9/QvwpNjwW+4l4LhwVTccMiUfO
zi0asvZegLgol48+7k3awtwTwDeSkB+vrgphi3gwqh2TA/hMehc6h8i99hHP3qmBIziPUqqi3XvR
IE/2s67DuVjCnk1WkYVclNihTpExaGEycmkVdPPhC0j05LIX0f+eBQmBDIqwJnwAXm/G5m1cWvUh
OS1elH9KPS+6w0N2RKFQkuqmyJuE7oHMcZryxwqNTKZNLlzTxbuNDmpvs5E5Ss2alLq3mMwKoJWG
4vQ+2IYWs0SUBgdLZUPV8sA9Dlge1Yf/B1bZKwk3brfbm/FCQXrSh1Bakd85twD/LqFHb1Iyw0bH
TC1gkRpJrdf1fCABMlaH4T1IUze1gRdVa5ETCaA0R9gfLW9HZ6CYfhC69gRjWmLv9dwaqoE6dPCG
4o1voKhuR6CggEx3YhKQDp1zn2UX6uU9NdSUjAYq1lxx4Yad+pTEvk4fSXAwexEbFKIvAgvBdYfC
NfBgdkFzbzxLBPunQEhNqI5Sh/N1B2e21yyH7CG8fFEd7zoF7pA/dE89KKQ6VUHWokM1vp7DPnGV
qKaZ5ocgD2rDaibm9lPu1+Qr0D0JeADFbVokkK05+aDWXKby+kW9RJEDpqbF7VVEw9VItPIKyY8m
WHbWUT2MCpFBWWaVbR/vkbK/HEddyxRaEpwJxMElVs7gwiS5UYYqxHGr5rzRX2MPrqK5nHNkvXrx
sm8lhjds38s6vznoKSpWuqcsJZeUlelYwQz9CHWMx/e0MusfNnWfmxT92x0OerprUbnxCVCO3J9z
mziBEP0U8sEZt8viu7I1qH5a7bnUuY8Z22qladgKgBzRp8AevIRJyAiSK/LwyFjVmVnojngD1L7g
z9PudvSESjJ5XFxWKPfwBTV98mLp20EK5usLvyBzqpTLWpozjJlYHDo85bFkR4MpV9mKUdLn2adp
TX3gqGrvpje5M4QV1J5pNJk5RMCVNVjMG32jRSMW7HkPHLYVa3WoXtdduDKXKKiJb5QkDaCSzzh/
lob4hNbrqsOHEaXJYoOZvBOZrcFPReVlyCErJg25u9ZsXejKyKT9suFsrwWEoAxH2E6w204HH7eH
OcQgV7nrMxJ0koMnKsxfpyaBvKA6vaEXdDF67HMzgtzrRJxrXQ7ODT05E8iUSrBxiP9ZIogWQMyX
Z5IQhCvBZgENwK/loaAQU7WoXhQdItRkU1Cnn0eU8zFTbrsw7j2ru4VVKsM2cGcJPbVETRoRz3GP
Ooiv//FvK33/gSAi/D9wPGRZcWOgU/YisyC3bCgp0C+aEgxLCtf6CMUV8ypA2UMLEQYx0N8ejJvf
ioQl1rS2TjW+Ik3PqCSSvfhuHCdwjpb3UJEoemlctJB9otATydY58XJln7bUvqectt5MjGz4b66l
raGkFVk+sKsKt2PkFt4E+Rh7GFIyqhPq/+wfQK04XaPYwv4aqbs/hdBNu2rAUtWfEMdZJZlWeGBG
tb+9vBVVM2wXiS97uwAPbKianqINmM7j79QUX3mADCzEsw1D2ULDJlUPGj/PT53GEGABd2YtHvAO
nkZGe6G7+krU/nx3orB4yKWsf5oEwC8I/Vbp9iuQHNzyujKFiumCc9LxfUmxnj4Je0f95qeScAqK
kMDGQRID5dfCFSzN+F9vnICFsE35yjyLkaM/i5bkHt7p4ROEn4sNDirykBX+p2ODEZc0bK9JCAuZ
FZms3oBCVyeuoPLvJAUbrnvPSWwjnUWxI4MYqVn3fZdgTL7Wi20TgV5Mv6jXj+80usnfjd12Qc+o
OnE5Fur7Q/f30JSDssRfWnltr+wrESuY0NH9BHmYAoAek81iKdlpH4o++rgR4RXEoqEB+rFi0tyQ
hx6duUTa0h6T6yCWNVmYyVZzFbN5+cMjRY8E/cRlKj0Fearr6jw8BXi8HVQmIa4C84r2io7O2OPh
PokrgEFUbUVtcPqbvdtcRd2fV08IWA6VgLefncJ8+CV6VPCtXDssSzUnDxb7Xj6NTQoOS8amrQ4u
RoDSgoPuX1tLZwIKgi9oX6iWo2A6GF3W8Lbwfk3rNRwfYJBvSrdoDNtf89VO59foi/M21T+nyrAx
mzUUvqANV9+e1GXEq0lrr7+PCNv3eRBz+oaCl37yfNQqAxv8q1vnvThEdAT0OnFprA5t1THH6xt5
julVFZw3+bjWG5xiQvOZINKcYnfFR+1r2VTBFcHekPffkt1VSzAfy/qG2CYzFYN/jT0LIy4+S7Zk
yni3y0l7zbEEYHsjbIhwv0mdDB88GIZwfju0SQzNp0/5N1KKs5GxJRr5oVxWYfygAotqH+uCxOZe
Z2ml5sGkOcnG16jF+2H/xGr4FKKyY2ZUdYc3y5WnHBk0WVeAvviw+WZ34X1tuJ1218GH9Fp1fSt+
coi8UTfyt4Z+JRZp05ceHP1gab5pBGwJZVHhka4CdxKfdj+59mgUTbiJnmXynzNqKf9E2Jcne8o2
gmO80l9J1zTRrFUEb5VYI+gm+JthrT1sZRONvxHbldK+4Gou9QxFybcscltC4tq/qCnO2eAyqxN2
h0nqEaHv1zzJZWS1qfqFHJ+EqBEgAR9lg0JCcD0O6/Am5GNY+QUzKS1ofG6UcEJ9ElHW5mYkMZWA
YrCyusR1XCEyd8FleQsrX2oioXr2/eVDwiFKHG0Y0zjgSpohHvlOkQXEo7q4cAOuHBvJAiEHx6UY
FFFJWTmMAL1gxs+XmOyN0cQOhZtkM9v2O+tKz8PQaxXbayUuqs4DrYVZwluZn6R3gx8tvSahlBmc
W+7iGcFp1U4xIcBeqNyviMVJCgoKLtP9jJ9pb88t6Pa4xtiUxP91+xQ1mXk7j1hOXNoEO3h75T6w
cwM6l+su6PUBcrqL59igS8ue2+FDnUAE+MEF1rLmkU+D0z4BTzv3agaKl/mfyJzpBfC+OwjVjv21
hh/qfFjOA9UjngGuOXIVwBdhhyqo47vNOAf49/dC+gCoEjizxP0/ZPBbHYiqpgra4KW9YnN1M2Jo
6brxyMLEAW1wIxfuHok+J1rVrKnKuzAiTwVff5HhawMTmCOuhRMZIrHrVseQEECTzQ4i0USw5H/v
YGW+xqXUu4OwR04+Vg1LrmIo77nBOUd8TpShlj0U5KetvsooCbuXdQlNzs7kwyB3/cW++actw++v
0lD/GO31WrIWctAskTrQybJCp2UQU88sVvlLTa/bX8cr0sEturxOBdbuEz3anmuleWUwLmqf36zj
Um2B4Tl5dSGdzVdmDSvXO48a/Qv9FNl3Ttf49KWce0WtpPwEcs43zE4xr+0nU8NzrTn6SLb3YXFi
Gk3Oo4LacY7nTuixJIWhr24/QcremJlPEBbyKp/cbyi8pbywdW/6bvZPqociMYvyCygd6jyQDSXj
JQcxAgDOrqAKIg4J0G6abIfNJQqCVMf/GcoIlnOXkWvttn0gl/ASeBDJboU/SRlOx1nOH5i9ObJ4
DD9Fx6zujdqrxiYVk1XGDHGhEobGbCjcIK72sjbAHqkm7NitdbBw1ess5hFd3/Wy2GjSGmAVBrXm
YcS3FZlhhbEvCrJLayxlhNav+P+G73mwAFHgDZvBuJGAjFlZ06vuCRZuCGOGcBClbhXFjLdHoY0r
DX7oVuwFUEU6Zbdkf0raLkOw+JoRxefoEmeSgFhR/XhUaV3vJ4NAsLY/wmAA4Vd9EMY1UkLGY2lD
DqcAs7yt/hne+HxGxsE7VndjXUGUnRLMNsCwYRW3bA7QZMo7CmW6+9m+qpixAYWmXKM1Goaan+8I
U4O5byLJg0sDR0DbE4m+0L90bskWK3R4Fo29dv5LjD86Re+qIX5ArRF4eESYKW7QeQl+Xi7E8MoQ
fONzFPmJ30U1DxbxE1zT24Ri8CShROCjkwxb06+xJA8JQRNEanWu/b+AOUEurScNiWzPMMoVajXi
Xkc4LmVJumr7uMSouHhq/K7Mn7f6rV8E5pxCVYCILPBWvmF9luee7ilmmBOVUwRHgLECyqy8g8Kq
Qfaelfzl3XKC5vzLf4rAJUq7lorzt/kJMRKbEJ7XT+5axfOSp+xX7QxSulpks/GRJ4RFJf7nbRsp
/9F+cadlY/7hmbS9QV0sX5X5LMyYB4Cmbd2Bh02nHhMyz21gGqR5zD1gtB51XgICLF0AdwmNbwEP
D9HMMOouhMidyW4s4B+d8Rr3cbvXJtrrspLzXHGAdv9QxCeGMxYme3RBVDOuFdA2G0BRMmaydLdn
IesCDjejV4Ge4qYT3HSi+q5uie9NS9mwtaAt7Xfw8JxSU1leTE+AMPjt1jIHd7SIuOd2h5dG4R7k
opO1GEbISm7AlX+1ZDiwoEjr5fC3ZJXUZFt0JDgblAM6jRPXFwxNOe5K75vLX6Qhgm8WYWgApdyU
QXiKQBMzZt0vsXmbOqPhczMyHT0HhJjEGridxHcr+JyQypW71qtqB9s7zAnXZXV7LudkrXcCBKNt
w6QcEDoLCNjd544gkwBRfkP6Kn68oP3wxbWdZeABUR4KpReEKIwfGXjWmSc/9zPSWMPMuw1vJTkQ
cIAabsMJOl7Jace9HA/hazkk+2Tcv1dXfDAw/sSUPjXPW8Gb8k+j2jHwB7dCF2C4rEJ6pndZfvH4
BoR+bynLcrFjqAoydydF+Q9NWI3bGEMI4ncAzpSCDQhjYMi26/n4wFfGY6nNuqyjl3CSdOYpgn4C
KnT92cEFq3R00kxWB87Qi7ZVpzS7B7UPZxJh81CX+ia1IK9qWc6pkLr3vUt6N5TdaiEr+ARBYH1S
ykN6dJgjgRUQ4kM6uzaSmec1HnkvTBj9YL+6JrZNFdcuKf85PKdGRtuQaLwvBX+mwT1SDdSzBC3t
AmCtR4HkqW7aoYMdeYT+ejYPTHlXgaKdd/1JazqbBCFcRDUq7M03KJDWg71tzhQDuqs6xrrdCPrZ
0pbEtNB7z2HMW0cZ8bc9fTQGwJcIXXMAf1G70Af/uJcVT+oTegP1Oaa2soAnXTGWLA+I0HgwoPo5
EXgGCbg/lMrpPec6bISqfa2TPy8U4oTsLdZzikfXqo7oOu/1ga1uhFKCBvaeWrYlA949VfRK03Nk
4WtujulxdHC/lLfjKF7zXXRZSBJqqZUQpFN8UIuQR3/QoxPpAWV993eaRmegVJfbuVXWhJ4cCO3K
SaaNI3neXm5hk1vr0FQX8ChiMVYF1ZU/fvieizI189p74IinsOVQf8LNuVm9Kx1FyCMNFxY0TiAd
KOf0+8TQyXlGwwh5WaodFaJmjYLSe1QAOynf/vkka1TrQilexd4QN/yEvrFl2bHaT44IDNPNwfNy
f26Kl6SmqfnDM6pV3IsIilVTrx/Txx99OrARsqQZ4X0Q61XGXtPWxdqCqbLSIFQ9vug1nEnDV5g2
JiZI85HpOhVGwk60qjRlBY3ih0XiY1vjqoWfri4jxlfcg4JIkCGFt5FIs/T/pMqcVsYz5NVVMcVL
DkoEvK5IOFopUb792xWaD6BJFz4F5NSlSOGiBGlmNdYhZFdM9aVNaQM26YdRuZb7PQw33L4Vi8/k
scEbIIrb/TCNkBEHxOb/+CjQLXmqNa9w8ZJYFY9YBvrPY1X4/p6qSf9W3S7CUkkDLUm1IKlTINo7
8bZu2Rrn/puJNGp569M7t4wp7m9Nm5ZtlxbA8ZruMJixV2CoBVv+qFois/lkHcA+EYbg1AP0dB+J
tTR+syDgpFAyxLVmsAW2/9/scj+Aof5vFysAZvYoXV3rjDTzcHmHdIgiStK9Rt50oZkn6Y+pQTQz
vJgNlWUx/3eMP7fER+xUSmEf17NT5TxhIXSgQt4ki6h0GUErZC3wPZiwfY43Nj5rrmjYpvJBMT7i
ZSTobzt/i6bgl6nBUym2G3ovMmH9vg5LbzsrJx4FHV4OayNAC+wZl1JhBBnvgosYlm+7yAZv8p3b
RxKXFCvVjQj9p3Kn4Yh9UNAyBl4Id/x0zx37pOUrH7XVZP8SRX8mvvIr3MMxojCq02lAvkFhWMEN
b/VNRzFYnSNs0rLRPoGGSJYdVy4QDWC6APijF6MXzrxIw/eOlQLNvuzeXLUS4y2seVZS/3bmNxKb
9iYjG9/o/3pjVK5G2UcbTQ739dqUIYpzkOdXauneCN2cOQxVBpGeFSX4Z8Xi6FlzujFvX2VzvoHa
kih1CXXqPSL4YSKkpACzGa217GaRh3nzkSQhjGjrYOrA1nvYHgMf/vi011qYiKEiSHmVF4SpPSI0
2dnkinHmZHrJ3p2iKWXXLmQdeGNhv/rWl2G3HE8PCjFTWJoXW+ybOz/Twxn+Y2/n5PyYJoik3VTu
nMX70Szeewex2eXFip0iA0lvxlhkw7gnrIJprPvIJ2D+62HiwTij5ekRqvxEsrZ+7PwDe8XLDZvr
flMQYZMJaKvtcvcFN+9hr/K4vke1FqzL78dT2DhtRdmBUHxqRKcqDOMZKKhmPOeqj4kDgzuo85N7
zyjlHo8B5NB7DKwwDMAD1hTlXlPE5atCQaQtxLkeanmXWaeHrHto/tUL1Irk0j4arzbGWBnURWKs
3UQt6QKQmncOjwMF+0VOI4tH8NGsl5Ex13VtRLsy2ma572J/JBrChlDeyer22eQGmRlTtcM5/GC6
fKDuGoL0RaaxVMyskQDra4I+Q4SyW68rCmxPxjIsfJpEFNplH7qaOyNxZY8L47L/uD8vW1Mmx9cC
lNdXLCN1FtkHAgyWdpuPVScMO4StBnN+ObhqbyXzQZO6pQounjb9QhXaCNRfbSqIkJdqppVU+JA7
EfeDc6vrc3gtWDJY/eSWBc87j/wz6468+o7EXVREKtBSXbhyy8FVTedr9L6xAlrg7aB2QocVKeb2
2Xlzk6za9d76eYLp6jGJP0Y4ssRbTPorzrfhSFEl1vKgIzFzmK5s8LTCuClInt5prGhX+8NpgDMu
mcmpwVe8zeB3/Ij3tUdfGZ/UabzPqgoRTmvINtdUAs51S66ux9c6kp5DifS8n6w7Jf86q123cVRn
IEHyZm7J0/39XkJAc77jCbemcYZ2Arm88Bo1R1LTF355xsByzu0CEbP6rce8zU47Vw6C8ZkerfrU
JUNjphLrR/CnQlvXj3pYrnBWabK0iSmRP+3yJoxXgPWKesiqIOeLgES5Qvfk51Pp2/8CXDtEAmJI
gKy6PF0MNTKcZ8WqCSnW5DMek54meaoOXU6L8olccSTFdToux1NDfKlg97qlurjlnNlg3n3RlyPr
TzPebtrS773ospZoStc4ZVS0zGF3suY+hbJUngSdx8keZ4xxahZG4V1K//RflClgccvzbxJyZ2gh
cjc4krIYc6AH3IKEl1GYJQPxl7tqbMH+5c6tKu+EQDEV5cYWs6V1N62bCq8jY6YTPxbvbQ5SrD7n
EDgcb9BZkxygiC9I7KQXzbmswJtOhoWGnAL8t4Izo9mAVOknVjSUeFUDNwj4NcHVSb/L2fbSFzLG
MubV9Ry699JEg5zLbO8xt3z2qBohcC4oQB9sMHB6YkfR19AEBQ6mCgQrokiI3CiAf6nyeYIyy2sI
lTdqvGZuc0p7YdzRc/jablpF93bKAOtGJgYwVy58gk14Co3WZ4KGw8PhJildwYz6fHY/ZXrJt9S6
r37ViAJyn/mKmfU3axezHgIVTbdjdRGZcfUSe04lDOo0vUTXorzi4gzYlBjhrWXLHrYTlrv8fnYF
7AdSpBJCiMHPqTOgDDaHFBFwQCurISg8IrSd+sFOH++hweqlVrXKnrrOon0sMIzj6STk2WuM56xO
AbWlqSO9PD3KA4C63YnJIJtOanrXJwWdRLbRhBQlbPom1uhXcXhDQ3eFMHuc5vhOdHyIkLmlI/lc
lSActAY3b0oMFT0vC1DUUHuZPQp6vqYYvIl7pLj4UdhcKubVkejl0WdEulvIi5mzP2lKBRSMbiNW
uY0NK6Q42OCKq20Sr0KZaROC0XLo0RHYwkv8g8a/lOLo27OxLbJID5hFC0eHvbqEzXH3azxeHRlH
JdtwpGkGZWPHGnuChLZ+pKOVgeTVkK3/21tQk692lq1YVptxc+gYoCSS6BdQBuzAEnAqMOS88+ik
9nRAYnf4sDP139Vp7O/UsIqVcT/kLzaab0IlCNRT3Iw/N0Nv4yVJiuQ/lBPDD7JkH8fncANGP9eV
xJcL7jScQucfynWK6R+APP1yyRyEEzZ/WT2KY5lkMRFJGXzuvOCAl5bOu48EmE3rH+2zKGDSrVKK
nZSAu/ydbwRNiZx+Iq26icohdDyj8EUWpiLfZgFqxaKAseskgtUyNog6FuTB3STNPADS8g/Sh9io
aBNZrnxUDR9MOKekzS5yiIP1DTb7lWsZ79K6Pg9JwV/MN27uQB2ZnGSVo0oiEGTKf9uvZY7OxavW
QCMT4gE+GBTIV6gEr0xlcZRtfALSm9qvE5jcRCRuHKDoaWdD4gjxcZTsf9T3dktVqd51C2xRYW1L
lSYMGlQSrKf1AI+JqwthodX3dKXhERmFuqYjTaWsXFAE/n8NT4fTBrYLEgVmMaUXkpkFgau/lW2+
fHvscCfo+vvNtWh6mFF18jhSrdeh5aHK8tZAzxvOLAZsGprOaKWK/eV+cExZUBlKVFSNQmk/bCMU
2aO8YTfzQTy0U9seh7NjKCLHTO7uvDmR90PZswbsHkzwDC91AAuYZRoLNi9b1IroR6k6Mp7ck/9O
HL60k0B/IniD48jkVsom/vQT2rQyYh7QzzNgDo1+t/6Zq4/1K2/8sQ9MNFUQdY2KCQMatjYffB0h
BIyqXXeWdGnLqdP/1gBDJjRPmOCCLz99MTwVi6ob9u5awAVnL7bdi+xwBwcYLgwerkuR8rTH795H
DeDrtS9UO1vdluPMAypYXEgEIPooFdMuBeC5I1dO4wbYm/nu+S9tkANPZ/afbAvPZf43yz0WjY4B
7vwEOulGfEgn/lpkg2KDCqDgc97HiTzMS5et05iFomqiRSU8DEFSrky6UizErKO2+4FwtdRYEyIF
TwQaE4aoeg36ZRP2dqYzDw+bT409kqy6tS3yV2YWetL77SNt82oNkCryeTplTvZiRsSlz0YMmXcx
id+hqWGQFXebKu/v534SaLg4lrbyxSvrEC3lR2h2OtC2cuX/OvVwVa6ubnlurFUWlUcEhcXgd6F7
6+IDF1RGe31QfngMYL7JMueMPbCEnEiOc7ZDsuCEw7Nxpz6jIGQRI5ViYGfsIbSr6aFWYhFjcxd5
OlpgZormXfFaljsZVss0xl9uYQkPWGevjeqgz/zbg6IT9Hv859R5/mQQR7pWX1uQuPNehPlNXw5e
tV1KOr+glP3EAQHW80a3YNKY+dYexbktk97xx0k4babm9oDegfRx84B0zkTYFMb9AIqMyIV9bd6P
NKrmnhytkIjmkScV6eV9SqjUqFpAalbPPpf+2uTwyx9M5nb9cdVNLizsU6jG9iNxPw7tKblYwpk0
OT2WCGwdSticVEX+IRIpli4I+6TTBkJIaOR0yuNnrYMwR4l1vQgKUWpWVkw5pEp87eIqD6lWT+cD
RaJEWH2aEvqsSi26uDXUFT0wXjkn2uPcEfZuFVe7XkO3kA33cnZC0xICenwOjKqj8m7FwWtA3EI3
LnJfQEORed+hI0rlRr6PKEBH6Nt9WDpxX8AvbXg5AxxEVcdhLs32fBDsJhe/imyAKqBnSwWSV5FN
joxdM+DOFMh/D2NlIkEqsiltebsACIi1bGRaysVyImBQVPNWd2RPwk/d7mWZC2PYZOUsJuykFTOA
kdNLWh9tL5LxxvWUtwBpUlOcpIVVWbf9rVU/xKFOY5O48vdBB21/IhNhakYmcO+MmoFf/KG/rv0D
Br8EiuWTNntI44D4Ku8ITI4stZVE+bUATZ6EtnWTaFj7Fuqb+3Y4o8LKqb6/NW+3xi9K0kTRAYIh
iEe2/5JL1U/85KdUwa7LdFknUhd77vgdT5fDKn8B9xgK6LNDmpNxEmZsTOfXqPSsEEFSC7hInS4b
5nQHMvOSCfpuuQW30Lz6iwW3jF6mDHST2GJnAJW8PA9J+o6bfw8reF2tws68iqziOrGBxA10lvn9
ex8rLauW+GkIjvd0CNmI4Yn9keZuvKJVzHqdLCHdVzacZKKX/JPIE7iiOgU08ILUEyUxcgnoyH5P
gZAgCiqSJ9f+NhogVujlCogTWertBa49YpnH1CbLw2AXQfYPzV7gAlKXU2/o3tX0gkqra0F4sDDn
2dyKg5cGEVhvGwiQcunc9pLDc7kMDa2yGot6BlEdJme03e7VLg1VQXflRzGg2BxI5Kxhl5a/7Gu8
u2tp+B2aTp14QOBCo1WDKygQY4rBZiuC4wkJpxPFba4t2DMNh5Ap1lxT1CUxZwb0tBhxZEi/4i0b
4X3xJlOUtKqruV+YATZddZBOBNPx0avnZQxcOUnbBuZIbOkBLJbdrV/JD7T4u3Ou/IQ0RbbERmEf
eLyOn0HlowbBPOJV5MnbGpptuNowCwUCaYbq++VfiWFjJ1kuzyZVJi5ZsTFBVP7DWpDjGtbpDR33
6DfX+KwjP7eZJbb7hSf/WSl0wH2l3ekPtE41QqfwVOW6xo3ONjUt5kTgdjlAQEeqSfm5jQEshBFQ
BOETPYemifhrTmdkuL7Ip378UCG0L7xhhKYDW8r8NlxMRy0YxcC9+GL0ui0G/ddo+p8+Ji0cwLXr
MnXH2qxaRdJToSO+ILoWyrAXsa5HUsg4WUIWyPCusvPpJwIqD2uOQc4N0mdL58EPHs3py0t1as89
N3dy8HpFnY+YtnEkZLNAFmJeuh6NrVjQe6KU7f8AOfANdNNXjG5Ia0bljJ5xg4I2ycMAVJnlzMwx
3t3qrjV/3r2J46bq/WUbwHD0qCJGDRvZIf+Hl8nRemWXO5Ko/783t2LA+Yr3spE4fBJXiPaaY48Y
gLFThZAG9GfFieGW/+sE3rOu4j6GJquDFnVp4FXsjkDLa6/INBfdNNZ4dHZFJY+H5YWKo86VLVMP
XtFjFF6qlOEu7BUgolawbNPTqEXAgNCarWKZtkOK+FEqoOWL2I2QIzPIEg7UnQa1iFLPlQpX14XX
eYHuF6WWwuj7dwduqnCmgNBUfYOqKNGFjY9IrLjq2tzENeUI1I/V2VwdRO42mXVvm4cwoaJNN+fL
bG2KuN1J3PvCg9xqDfBpQxxRwsEhK3PoRjsq0FC4GhxJW6I6VbobZPSttmjMXX1ub6K4Uhoh741n
AAjJ8zMK3wcTeX2kQ8dvMNLNxDouiGr50yzpAA1kQnj39t86p7eZyFOcu+lvdGIlbKFFFRp6BNoU
JMujV4ZMc0RLmd/5lGm7N2n/2mlH6nGR1pGRJoZ87/hxpedGYtBUtZjKCDk9jLMqVY1qrl3sBFG7
8MWWBs6Fguk+Qbpi7Mfn2/QQZPcXeYUiim0G+f071QnKV1yc3VTf6OafJ5IeA06m1MqgIYTwWxK2
87xqJeLzhHbwIhnrALwjNIeKsf8J8rHrZtdhkZ/iVes9nrr6xstsBhYqiP/9bys3o4ZsZo2+Qf+4
9UXQM5M/JTljNleFXx09LekTKaC9teUDYS5IJFj63zeqHuk9Cn9/o1Ykx7UxrgykXLZ2iuAG+4yi
7rFsGzT0RHZQdXtVovUNBSsnWlIws7WXyOP42HTc5ppoFlZhq/1gdri/3ZhqGTbMhL+wZVi/e5wT
LzNd5G3oGWv29Jg28dRIoQI0UizBGI3zX99WOoXyrx6QKKhgQoO/syFis/9Ohx4Z8Q+HTTbEwkod
XRFmGxR3pyrVZSZjQBR65o5luFC5JKFZH9Xv9sfwim/7Y0hyEihs4Py3mAD2P3kU0vCY3LE9MVrW
rhwNpXwO4A/t5TWt1vJpeCfhsBOYia1+aYEfJEJqDWyX2i4WIdIurgKVZB0GKGWQRGiUkplf5mi6
K1FgZeB5IcQNxNm7l23h1ydSheCAc8xc7eMUo2sJYr8yWh+5ncRmvNcB/R76nFj53fDKNvqtoN/A
5JGSJsnUuGrvLjrzDXnWurNtoboGdYPuFmXL+TpRaQedevY/oIhB+RWvd5m5THYGb4ZNvxHc6t3e
pTzZK6xax4Y9mIvrGxHek1fYK68Xx+qiXxO2LTXSPIW2hQMb3hA2Oovmu55KdteAdI9o7vuVRhpr
2mGIr2pnMNUhnQK+mNu1tZ3irz8zTJi0eGxsKiFCs0ybrn37PwDVvXB86NutoRRVUO6uuj4b0sa6
uE4hLTdiX9k6ulZqB7WL2OxY7YMt71OXCAsXghtR5GmF8pjfvGqj1p69G1LWL0nxeLnKiINruglE
pG9jyV4bBuj5MR3vbJNhBwEWA+h/NuJZZIC8cX3LfxPmm2SADfuXg0ArkbvivcHrxk2sAd3OqRHE
1Wt6koqUaCnncNLaK3WNL6j0qdxlutEFMOgy+4QnhgB6iKsBsSE1dQZ3WOqVM5u919AoC4ld9aau
uGByhkoRK9JDwEBvEbESKBIbCeU5E+oDWqaAFJ2KFgvVmQGWRoPHDOhcQx69YjqYTiUdvHGdmAUH
LRN86iD/eEhs/UP8wNhmtIPE6NWckHJrzwsZA1629wAVq4eyhh35ZLl7bhAIX685X4HFfmbbDkCG
H494KhTN2OM1lRWfNX2+q8QC+t0s/70ej2Ff98X2I3bWrs9vLXnZVsJBTI23rEJEZcYmAbpzs1Yw
IFAhAkS6AJ1ifK5GBWXMdgTNwkmFicEDaTwoPi1P5mSaPEPIwWWpXlbcTGDBfQuFg1vz1KRjDSEx
oAFFjpOLYVJWKEzOSvb7fTNaE20R1g4ZrwQhWwzx82XS5bsWuZIKr0uilPWsEA79gBmYpk83TM0n
Dm1SO8gyMteojURbWEo//iG4oLAsn/u1wYahQMyYS1f5O/cex8nfYJFSTb/BmZEKOTqhEBH5SFBm
2+IQxr5CuuLACi/oWakrg9AxrOf1/yQl+GmmMB3vV537ruI5wPhBS9seHsL3bekOX2/Vw3DJ46aU
MQWWB5ILS17qDWGYvZ40YV30FAsQjSQ86P6zHybubHXLwAcG7N3PUdVtqrwIFz9XEjoVOqnfH1r1
2EAweZ1Smwb1byLdW8fc3o2hFsGP+5HfW2CQZ+gGXgXWZ2Wbk+87vHjb8SuWZt7b2IaoPVj+2pxx
Zf8qs/WarQpgmkGLZpG+bT8QsboZm/kyfws0TjjqEDKkzkPhC8w+Z+xSfl9pieo6M8B8uEFYfl3f
oHdDic5hCThrf1NQc/rO3JiLKP+DWP9iIxTZkyQrZgo+3ivyB3utUfd5rxekfmbKFlbai9viZfa3
oEycwqeKENoeNpym6ddYfb8Df3lrcZKHbQBrWpRtacv6jb32UGJ2iXZ18yzqFlCe4PN8/eBVG3GO
SNo923iF/oyukyqf/QkcEQg3jLShDhbjEM9k5Giq5AEfYseq82vHrCepWSxs/WwCzgbD4Wm3DF0Y
iT2EOCIw4XM4T4NCgX8c8EpYS8kqAF9XRmKqymIXo56x8NBlFAAPiO06nsNdxmSwM0+IYjtLUYpO
VCqxvyFLITlAkZKnK3mSUsWTm95PVq0I4knrIkc5taMnq2WHGHi8ukPNTIvbvgV1t7FOudtqur3A
S3GZc4/TYNsDjF7q5sKR6yP2tKp23p6q1qKHXUvG5IhC6Hyf8ZFm4BnugCRW1apQ8gXR16S6FO+T
WUeCU76IUEH0RtqP/yJZ9bucN4Mb7TzmT+7wdVow5sMRV0ap7/IlHzN/gd5o05hk6Dn9DJL2QNP5
HPHI5wsTGs4IBYvLYZGxfnpi1MzfhFd2YYmTfYbj8gWGRCPmT3Swl8SWV60g5QQB1MIWMA+HJCjA
ZVzy1hOaHU6CW4QQhWWLaH7QjGLiTGQUkoskV3e/307Xo+KtwaYQMpZm85VNT7PQXIwizuvSTQ4Y
ipFfmKSTsn34VmUI8g79rrMwr40RWSqivL+34vIg/+SYJWJDYSZyzXzIYs4Ev84tl3L8+l/xtRV0
BpRm78aijibxF83dA3IseqFJQVbtMhDrwrPmwAG9O6KhjyNWf2dP/RSjyeQ/ssH9vFgv+Jf7lxsg
FmGTUJQ0feDGexZ0AUmQbI2G4Jz2/weLYZcj97m7kczVmvUbUYbaG7fWmojSHieGJn8ubJmpsEcA
nkCyS4C4sUDjCZhOI1+F1riWl7ifO77G8x0GhiYyw/AaDgvTwf5N5zwvMfdZIzTlIBtwj3YmybxS
SrvHdppHwsQhHV9XGKFdoMGsKbMNxPPV+9gX/8rdgPuTje0qFYLlB2ViXKxn0knYvqeOuZeWgawY
joNoFukmHgK6jRd7b5LK5CqZfp6IuPhX5ptEgA7DtSUlj23zfAhIAWrBDFB/XvUkjwRS0+GeU3Nn
SEesK2VtcaHPaVrUkLQAt30y2y1iqAhZstO44311F6DOkMcjr/5+EdA5KJ/WhtGsxL0u3KetRRpa
bIHbNKxxyynXFCgSR3zSQXbfiWyv+mvYYmo0A1Dr/q+nBcE9OqG8dX9cLzAGqKMOG6nuxfW9+uRX
8VbouDR84qBLUpEDunQ7ah9CtdXq8h85xxbIiYFqQG4SYFwU69AZ9uWhyjKBtYPfaYJLh1FDeQki
iJtm/65tMjnJ0aZ12l2aX9zBGtpccAh6OUtUFaKJEfCq/alpR0PUEXFxODBU2cgPAxvqhPFGviFA
AVt6V8u+lsraQoHg9wT9Kuj9SwSUcEryA5Ei6ZciNFxK23VHV5tBkaEp6RKYXjt2uWSiXA2MPEKJ
Q2whmoO6WhIvEiZYAja95WOqMuKs3+cREo26Gpjh07MwESLFAyl5iibXRZIe0VLcfDIbABU7fSgp
pUBpEfhBy6qS51ksLCpQtcu0Jvuw0UW8klp1wZ8g+JxumyPcLAIlmCXYm3+eqZ6V2s+2X45jfG5O
tjvhh+1GFvneTcUYCjDkan7D0XGjm4qYEkRGR+IlQjw2pRdKWmHSGpfoB8WBv4KOVIUKEBoYKNfh
1FyD7TuVvpuWMXkd6pNT5bgcwHnesYfKW2bF2tuZEZ2bqBxm3ucjAjzRZUtIaKZaTjT16mH0ap+l
7JUBYWT2cz7iMlSkq3FrAFky988RHbvYJBGUz5VlSLmwhxFG3HfbT5hkQxtnzokAvoZvB9WpAQV9
1c2pulubYVSPfFK6mAuwUV6h6P2oHTJsJzwEcF0WYPkbAPmqRJPLMxp8HyUy7B3fMWf6hjgw0yUh
23L0QJKjzlbR4F2Ewoz7aSXDh5AOlGbVtCXyupj3PPMFk0XDH3xa2Nz4bbkfcI6AoOt5a2X2Drwt
6qsGUfQ6Xz+13DunGBvrTg1f188xJYB9Tzuxmjc/4Z17Zm5gLYNa9oIGrWP5nJe3Bzu/Nf/ZxAfZ
z706IMH9Na3lF34kJmmQRLrKM3fjtwsZdDMn8gLLohySAUJyb8GmYNaaEtqaP8luxN3rlcbQVVFW
kNwL7Icp3KZwajoljo2esshKG+gPIQZEva59Hc89xTJ3FrMAEIpWu4aAQVBIcrginXwGXO9XUtl6
/P0aeTt72CY28nABkUDBuqg3McdtCB9seWKacw8zACTZ/1qAd3bW18YXXAY+eGb0SbWE2IucPc56
s9OhDstfSLyvlXvRK6Q+HYVu6Vb38KW77MSjttOszW/+DZZDmmi1puxo+MhvTGvb+D3wJ0zrUC6J
TfLmw+V0C1GnRz1yvmO9KDNEAPFW5gTWGzrUXUrKFD7E6IUhtzPHwo8suitDu41Ijxs53/Tt5ZpU
OsV2Hh+UZxmAceyjBjEYsJtdOOLnphPtOD1CJd/91KEqKpB+zK/WKLxCGOUDu2Hdvu1XfDnSuYjO
odASpvcu8ILIDtNI43rA72ZKbH0kudaC/uRIRtHdNT1VrhfTNwVSXniz6bfbpbowqbECLTHqsW+R
vsw7GZ0LLVt1KP2q/DbBzQ5zsNXAkT/R9wL8fbpmDk4LJ4rGnwDHRUsClhZKjG087by9NCJE+gkA
oDIWYRn1XOdR/hk9Qw/mgD/8mNYl7HtTlI24FmV+5klVcfVlfYc9Ir7uZxO819C4QfWowbs03LEn
6TgbBucP5WEte0af1HWazLdhvfGJkswiRIIm/FUy+KstHV6kx2TFJrg8WHlocFDNiFkZdV6HVkUo
2ppyQ9ix3kB/9GxUsiI8JqeJwADUpnwXcCHwyctmeTdaQ2Frzv4YAiP/cSurYOaQJSIcefv/dohH
luSeEj/D6c0eUZatqDgn5PIdrqmW+RCV+laXejPX3xY7u7FdUJX9g2MKn5TzD5mR+FKKxz+sSmV/
b6bB2T3i1DNbgquzkmELGRtedWb3EnQoQb1tRa0DT7NsJoZ1tg6cm7ttVK6el19OO/ZDcxecUW91
2m73WV5GbiibvbvKumQ6yho+ZglI3kPKvpZyVe/NDRtiiFc/gmQiI1E/WsUAEWQIQ2zCdjgE5yTA
qb8iFYfsN2cVdzVa2mDvLr8R5XDr58s0LYR52tquSXLGqNUSWnFaQ8NGzoKWZ6Ibs41aY0jCyZ81
aFbBxOBr1qfokKhOH55gegJ0Oya5igslc58BmFKOHaf4MPfKMP08Ryt6vNdrGz98+q2Avdi0D5qC
1qA8SW5nQyGetTXct4G1V1CzXaaoxU3qPkamWHvAM2k8/b4bJWE6uP9i4FuCFqoIJlcrJ7G1AAGG
9q6IpumPDH0Z6PWOlLNd302jPdCkT37y2ByKGjeV6payxUHg3ilt2ztCWsQ7ReL/8ma+ziHt3IkN
1+zNhNLqWmBU1ZdCywaFmAxsAhHnAPUq+y1psUzsQUiTIVRzL3RIFEX3wg7RkuyS+0zL0dxK3lHB
i7uc4XAZD5j2aQSBfjjVsoMx63R6cytWUylBZl6JZhdpOTL+plHs0xdGQlZtBznG3do5x10ndnmf
GqqhgOrkJVYTtd2w8CmkeEmePC/L4mDvaQJEb2GwBMwYAqVnjSEtnYLycmbOd0RHGk7bRaZ0zIZe
IzVMcQ79XBRK6lyFs87yQBl/RK2v4JJjYrsD3F4Mf3H+7/ZJTCR+M5ddofBZo1lddH2FbJSZIdQ4
QSk6Guz6EjaCNCWhfhs45A3gG4VjKnOTGRXzVGch6flopsrOXml9z72qqzmp34CGW30CfpRI4h6o
WyRrZY8LMmzbaoJ7yod/DwJX1CQsAuXYldB8a5wRwjWbkYnW7siTau51Lz6wzXixkNb3BYBa5CvS
xw43T5JUWXSt4PT27Y2PLN8zXAy8fD8YSRjdo78LwB45Au8GZLgrNEnzGGwg/HuqO22hmrtKutoD
X0tMalHPGbpA9iPwCqctKZ/VnHd8Q8INoDVyCdiTxBLx13krqZ1xL/E2bELs198MzWdtUkCgCSTO
C8ta9zxW04F92GBReQHDh6fGELaJd4syPNalQ8+YNetieiJrhDQJL8x5SiXSpWi2f7ACikEzXRoI
5tFi1c5dFl0qQhMQZL34vZdiaOR+mkzzYc+Dfcc9OHePP9QH3oJxP+T0RUw1fvSsn5sKN8fjv5zD
GwBLSY5knJv7aXZm2TGzEh3vv4ZlXJMFRebA5OL5htXWXu9qf/Q198SFZwKjkfCG3ZBZ7LRF7YtI
4CZPixQAIOBfAAcmwpCzez8OMSaurdPQ+GFlQ8vWFAZiYZEjjFAMlANqX9PHWxWyBSAeH9Y7UF3z
XXCMRhfwQsUh7nxGF1Yk7HKBh/evtF+l/zo5Ay5jhbFPeYg06lTFlqeLXkpoA9tTa/4DP8hzBlRW
B9PUciBSBc/vZaf7TBUxdCV835BjPF8LooyBhLrdZTxAtW9DhMl3cHJB/eM1JHuWfQUI+Vvfr1oM
O5cYT4bqUmUKT8Zr+DoCNwHXW7XHwdc3fXgXQr5b3OvcKwG/xtVaeP1qobGW9NiijKh9cYwjlCi/
FLdC0F5I5hyJXn9OEo4kgvqM7++qwbAfFUOWmHS/pJ1KLDuwjXRxyi6xOCIF4rrpExWfrDPBYNBj
DeUkL3mij9LxPa22xSR4Zaz6DMP3CuEfhrH52oSFDZC/20BDRKijiwueeuxP5+dlYx+jxcLnOJJo
O7pD9WVPnpRsK7+OZ7ejMN5hiKOtAFcjvKrbpr6q64laJaFGlQZtPExmKyCRmS6yPAGAt+1fhrnl
o66XZi6kahUlg6nWiayPJvDmC0vxpTKeps56cfp6zEQPvenV8DMfvE6rAFbArl3f0G8FX3fN03Nj
cmpiSS6gKrvll+Vwp3U7V339pFBuMdW6xRLFLoIz98QVo8sUxoXGh2l9aIcT6GL9Hi6F/+VZwPKj
ECh7hbCwHb1rHvhu+qd22GMo9Ou7Lm5RZl7TGyvWhtUKW3GHWhYGUMaeFLzy3SQgTRZKzMUl62+I
ljlyCZmXQkEjicNAqtpbU4VxFVnCAVmcKmMvXGRFS5/Yjxv42VkrbjoV0jBicpDAOvjoF1ugvDDj
QSe3gxENNa07om5vwDZrI29OGOGyNPTUNZpqEJzxPiYO8aenakyH8u6jodn4UrcK0DKjb37KKebV
1vLmW6ljmNsujmcv+YPCS095E11lHrL996rGrT39uZKvhBNoz7Z7RXDry47jwPisYxf50BkOpf9L
VwEJd3R5HUq69rrYMUDmqakemCrofqSF81WHohQ1KF9ukJ5e5nzcnlaoFFadZBLyeRj+3j188VLR
czQzDDHu4keJ5sbzfoPJKtGkhran1fFJY6gnrNzxW1luVMYh3UbOLXnCVIjB6FYi4czHt/c8/MsR
n5hJdltiLfhoERp2D/xGeW4WBbiBZ2ZEdvI6h8nSSC6n5V6TYtDD1VJt1RGz1JGU7DGusgOaBPDh
A9ZPvHqFjMIK3Ust7gYfoscU/mP++q/Exfb1Zqq784eZ6LUcdoZf9UfsMEufwDZ3Y8nwZghQ5wfJ
v5sSsPog8LexDpDCD4EXD4PB5EXr7QLR1HXuwbltGcgfwTmDrSZVmNOLa61upYcXyC/kBHicIuOK
ZOrxxg18Uu8+GRW0zo+ptV7AWAuNpyi2Ta5dM24NfNhRbZ7zZagSdrIRZfXJXyHE3/1xypDXK94X
bz/VQiR938hhPwLLdYEHPf48Zkc87k9CmqSR3JBmYKf1zh5uBWJkKBBt/tnfJQpTWdSAj3h9J6KV
82ytPyODBfA7taDNMSeMZ76ST2zr3u1XnOs/gHsjZk1wchRGqbg9DqqgUn6klW6e4LBTqZ7ZOkzU
mDIyIUO6HNmzV509SIPJsR0otjua7Jl2HgFJXVpKWjHpSkuyYg7bZUxyEdRxYTXzDMJzthJUbUiL
WBpYjsDv1r9gC3rtRoyrTpPbLpa7Z7UB9tvUMjBhKsTSmK4MkDH8fMGBv/opc5PCiiW5E/MZCRTP
7KqNMVQyxogjqKNo/5LolGAlJIPl4Rr450lY6GzhSNfqqWdymMa2P8kM7jBspmadEIMbPdHxp2jJ
aetVe6giqGxchVU6C1LeviW1sVDLU8VoeIbSPftOVM1GprhKQ/kqVuaCiZlcZ7feCMWc4Hq7+RxB
xNNqfNdFPzY+veoGMcY306WGIbIKHInVDfkvno9HM2gJMbPkfgsI3WmBjNgJF8EBm3a8sDfI4cyb
fc2Axudlngj3wDru8CQvdnpOHBeJF+1d8+7sl5eUB8EkHVTeek03ta1zK59Ew9plqJxxpIvKj/p2
w5kfv9P7HUHgXFP8UJ8A/Ggxgo8o9vRWC+5y8Gzfj5sb3r+H8Pe374n6WnFhzsy/J4D35Ro7BC51
1+mDU+kSq2RS2PgQwN6ohkOpQ39MPUwwFFLkiF22ddT1+wcBTSn13Lh682Cm5DfVZqMjzbbs35hl
wqeGq0/dzW/SC+RWJgCN+fo0cZuMX0HXxvw1w24Z0BzpGqlNOG7wvcRA/AHn/nPw0mir3a0yT3R5
rywkKCPeKcKqRHOrau4oMx56yNIbC+W58bXxitjpIAJ+/mqPCb5S1sau7p/HZCPDYpijtKIACOJO
ky3hczHMKX7z2XZGxWaw8n0o+etpKIHMhZcegusIDkaREGp4C9USRE4ThjFhEa61429Y8Wo3Sxqk
VPUYD0Qe2E9yOWoIeeey9UxDCydj5KJxEym1sdSW3zF61oDNFEJ0ZxwXp/P7D7OolTDEIIghxvhU
O34jkN2rsf8RWq6w6DBdYi2IYbQ/06A+B6D+Isjz+dZzozyflJSo+ko2k8nTjrdPOwvAZHOfUdYJ
2hJCkgYde/CaM4HTujD1/8k1bGVXmTEfMdIoj8fxI27m2LvpBb/Qi6Hwvv4db1yi4vHMTcn4mdsm
ML89dkgry01T25B/z0wSW41csycUktlLSSSDVeocaHu3dFoPANtB+/vXjNVLg45EDubfte7hEjmk
2H41Q/iN5fgctpxu1HPBd8eug4GSDy9JGkEbXssBMR4XnVKi8cSyMaCgQFisJthDWbjFYmbdy5O5
xujeO8igN8qi5LPEYt9fNWiR+ASDq+8O92pH1KfZ/SMoImLbBpz2lhG6mE7vFzaaAza6FukYKrRz
5QYFlUT0NrUg3CkHVngePRu1K2llD6RORxUbIpqMkpAXMxgx08BPPq1dxDZ22TBt3SfbvYda7ECP
RJ1VDi5szFlpb95FtV27SdxYC8XBJ59VncUNrPV/mGo3AFvktjb9XhFHNvdVwUFe+wUzGWoN7hRo
eHNp6Vtplo9uuzGElnvA8ruNzY4jlquHW5c2LOxzSYOq7MrNlp3a7PsK/2HK8B05JC5WLLbuQ4ur
6VguIJetsvHyLRAnPFYKAd4R3aOK6x/8YGnukJNBoX78U6R4ROHG33S82wQCRxhHwU59DnuVB96J
VCxwqgGU4b9yQ50ucuox5OFvUFC7C9gi5Kcf1iG8V31qYscStE20EQCNpbCN8TqxHqHn3i3SYJn9
+aflwBoNYUzMT3EJDjzZBuxRKClO3LimBLN8O9a1/gLD8RgqoJB/IKbHKkCZJG02rWaApwDkiLoJ
I24lIQOjp4loXwbziTUWDyoq0ygMmwp7X3otyTT+3fQlOZhMd5kveq5MJR4tiDHzY6OJieXqY0yX
Ywz4TnTWdIgdV9+ozyNt2LxuC0/+xwq2vSnKM4523LhGGh5Maf3A33BQgobUEVHFN6Oz2dSeDYPF
lENs0DhWcxehOea/buT6QWbI/OE0UVNCz8m8ZxRv4AzwOptfSSvajjguknUJe/guiV6pFrRrZQDp
afqymCJ3cGfytdGcIk+U8Q4oWWEVS4AWUCUDUyl88QBKLWcThpe4meP/n9WoSoy9qzgYzFFLLV3L
hvd3Vd1fTSBI141zH0hz/IYvS5YZxMOE3KGAHCJFdB77OTLjq+3UwuK/MmclVAUYR8jU4YHOU2r/
4GJ7ftRsnmiMHU7g3oES9t7KYM0WAB+eRiLAkI7wmLH3N6SW/Rd4qDXiYgf+YKmL8PeotZPld/RS
co3X1kZKOHBjYYiiPjnqCLUJxpkmfUn0iV7MJpS/H42X9RI21RefTXt9LJw+4hZKRJDDnHARBLc3
jdxFm38ltgyE5XZ2MEH3YomAF4fxoUmWwo7K8VOGoTIuliER+Se+qErcozMg3SQXWSCNnnYh/feA
B2g5tZ5ICzq/2Jf6Zq+lQ38NGLMurTcD4m6XIK+NWxPVHDsrRVwq33Gfub+LG7nhsrTM9HFz9Q5t
X1mRo7zdCESwhZhaYR1rHO0gybi9+LQTRF8Az/Ptxx8mc1bAYPYjpshZoNpjk3HNIyU4jxKSZ/Rx
Gs0g1d8g99LGAUQMwuMB5nqJ8hJ0GAvAUsHXFRdGPbZ+ycTOhEa+MExU15P++QcIp5N2J3kW8ZMa
5bLK9+MzJYJXm1Ud4Pl8Iae+9BkQs76KbTZCwTLVU1UkliaClQBQw2hQ7T1w2yTgU3yCRDl1XkwT
ryoxEvffrqV/QHlPdqNclbTkSF/aTl19+gxAW6tBPjKQ90o+9zUqsuDHiEnr2OY82bA/iSirXH4e
tqlrGmnEgXQQ4Je88dNPXhXDyEAYj4IMcJDGXchQAN4nwHOMeo8RA1MuHzSwuWqKtJ3Iu7ljsaeK
pO7Htym0U8tfdvHhpe5fzGbotU5B44+wJ0WJ5uu3CVoVcdhl5Sve5fyDSmSjYrPHkBT3n7eJ0QQL
iQsv8Hd6Ufxgt7pmEAkwv7lwrVEwewzD2vq1MbK5RtYqbQ1zxMjYN6uVtScYtPmn4oyvZR2ItQjC
0tppK6kOM+1G9u5tgRKGyVmOHyXNmIU/7j07QYgLB0qdC/uaNaPLiYvh7JkueJ5Bz9uLXt25MBmO
ilF7qTscdqBMmUiq8ib/r0dMW6WUNOheqiVEiDvfK2YLlc9da8l5WndYjmWx42jAXkC+DJN5w8cg
El6/y2d7VHG4rtyRcvKJh6K3GYZAkUwwj4Bsq6W7j7GBb/J0tEvJq0INDQA9wd6ndVGmLyxImDiQ
uIQfO0VleT+rV/gFwAhEQ6ELErcFlp0m+MRKiwXHkuqL2JjtZ5ZcAunDlPm1h5okEmauCOTfwqrS
EEgI9026oZCzpcYaiLopu5EWbsuJavESetm93a5SF1Fta+TFx//rOiUlpbxZhLtyX+NnPs46QsXM
8bd1+6sQgvJkk/52Yp5KBZXjZdJY94Yc/jhnTjg7WiDDRZn59zOGR/BaePnd+jA/sgp4sFBjohj1
Ns9MVdzjD2fIGYZVNmTDXkQLA3iKjDfTS27ItRQGoeq7bVpk2d2/Irfisysm+9KCQOue1W3yI9Ms
v+WgV92AJr1tLLs5sJVdnKrxW510LDRzw/PruwKK1Dd/MbOzhDDj2AXKwMX0PL2CqEquf7mHJdVx
IN1kXoG5V/iA7ifo90tcrgBjXHpWTIeh2wTydH8JKSBBMFEy9+Yit4ayKTPFphd5aVEFGVlsXhxK
rXkzIvAKZdlhcRDmHTNpwHDtq/w8J3NvzjX5hvAzi29muAavnyfSg6emtOBX4OwBn5zy0UFTLJSS
huiJPP1AHKm7A+wBqM2/UclTEerBdBG5BaPSpatu70amZveJrag+i/qNBcr33d8R94A3P0OaP2hM
HGeWtd/imkXHdQRXbn2lcH0lWyOc8iK/H2FM2jXN8u6/RLa/iu6Q6AZe6x6BOX6ACqmbW6Q+6R+q
bPj7o4U1Ya0LED7js1zD5ToNxFhEbcXv7Hh9FjdIy0QKjB5tldUWNqCNCWWhhe5N52J0XW9sRC8m
fd2RPPGlnoT+JnEXQSerxbyUA6gydSYXD4P7JpyFuKzkrV1ux3v7qX2QOxhn+de3VtcJ1n4pVk1g
tt4zFOEsN7MQ8mZwhe/clE4QvYtLnCt0EOACDTHkJGZU5rEC49TL3vpHkT/AtLtKg/ImTjpGp/JC
kmq5IQhrPKz7Bk0ZNkgdM/qoz6prNIW/O543DgkWzkYDbEAQ3cpEY/N9TgW2w43+jtKMH2cuizrl
GYhrFrLk46tz88o39/T3E6zmlKxt+5Xp2mNzRwxKHvCTgE+qgOvZw6wjrRBQ9/JQnH3kmZphAgMS
vOKXi4jaiUZxd1JrsacIgHi6bSl8U8cP7iL2WHRzIQmtRBfOv0oGh23yJjtJEf8stUhuVUx3R+Sv
44XyrUZB0vdnzODMdOsWoMu5aLi5lUdTWaSoUAoU5YG/doqMTrkAFmiazwlLt3RF4ey76ni+uuUP
rsOqiJl2s8Qat7t4/M70dwFZQHJL1IOVmAQnbVgpPn4vLs8Pp3Z5090pnFGI282mWJ0xFRsm9b60
YABFAuBKfFyPoWwxn+hGjaBKDIag4CVLWVwzkxdD3b6QVY2ksBBmoDsRJE09cvDvKeKSCRC9ABwI
zoI1Q82ItVh+pK5ogxdhH6B2qlRS7feQGzQfBxgQRncTsVFW1GjLQBm+zJb78Wk2uNVI+305OLB9
rCPOIsovAOp66zBlZtFAtp8/m6sEO0JzFiA9C3XBXfyKhKeNgl3YcwcIVsKXqt1h7/ZtNRC/ctw/
lbVupXNtn9UxygjQ7o7PUfJUuaEglANNPGHnLnfBNFoqJoNfgh7uxgfdRz+HERTxmFb5YE9lEN8a
bVuZ3KPmeh60mQAEC/84WivSuJ+ND8zIku0iPNxtsXd+cbNpFhfSm/G2Jlca+N8ZRc1IJ2yN6aGo
mEOh7LjHhWGtYpfdzmaPK8RjKFI3ZuP43YZ/gO6IlLdVNii4toCxjHFhX8hIK6oQ6gBpu5UyIc/0
e8OvFfDLSG5hGyp72m9OSb0TQKJ2xvlMpgZmGdcCABdKX6AVB7toQEGihSM5WlRM8KmQ8lCSNZcc
KwwVbaYBsIZ0CdtjcBz5GCm0rXCRDxDjdQsOqdl1RF0AulIXhGaRe0anVrmMhRN8by4LVXZ6yQKC
/EmooGRTgu5dvI1SB/0OKz3Wu7I4SPCZ+BFupU/eXZcXZg1TbaRzUpg/lrK7/OHnQWadY3WEtKBd
SD1x+vs2x1uwVf8Bx7miLz19KjBNzw5bpq2L9rYg3t1OZWcdrlI9enHwstAUNIGMuHBLZsikAruz
HP+I/leZKQJ6X8znYPnS7tv7ACto69f3lodCxGJa3rAv034jFZo5Nn2fn/EDGwE3YED/oxy8Ub/c
g5rULvHW713TaMSoI7VqmlYOp0phtmK8IgBf4VptLRkUyDYu0QSO7GybeOY36MvBkz5J8V91Z7cd
CSUdiPljraSCCJJdQ72cjds2DUt7YN1CcC7hOkw9bPSB3PKPJHIz70Vkxa7Ara0QMwl7YhH9NL32
YXBhO0E/hYQYbQDYdAMZ76bdJJYhQIYzaDOWpBReqbqBuFsbta0OyTenrVXH7QofkoWoWBwnWk97
2ywuANXKlyBWM/Fo8yRMdz8HbQSxKFw8bW11OzYIHb0y358k+CCQxt8JT6sIxaZMNcX9lGMZSmLS
PKa5+ch6t3upsboF66gQKdaYZ8AtU+tyw02Pgy6aY18q9yjM2Cry2JzFeD06EuKy7MjS67MYe9Jk
SzyiFqNMbHneGFB4wYsnT9rePmkSJrF+l8QxApyssbqvpByJsZTlwoJhRwqj9yBtsljx68VDn9sY
km50tp+ESKExhCjoHjveFP1FA+qPr2vv65rEbqbbLL0V2WomyZICg6bZ8gtwXQzekTo+uPKgWD3k
P681WzjLbrvIUzl2h1AqymVYapIHZfNhlkKkO4WnmD+U3/iXKPsnLRQSVvMtYfN9rT4T8s6zxOLQ
xE/R0k+MIFmx4zu1NSl/B7tQmMoq0G+dSYOHjuSc3iHZoHdcSbMyjYdaZOzeWFcstPmzd9QBaEGC
+bamI67q9hQPMKVoYUeg48dhr0IQAGJ3PlkHBKyE/2UQqd3hsE9ubYfKie4R0gNfJssxBWlINRol
gtZfLWsLNFKKg4CTEQhSD9/Kd0g/h2E2zA+gMGbrZ9CUPs9q3MisVJ3XE7vYL+zu92CqZ+lsXXJd
KgKjD88Y/mDnGT2FIw9TvFBKB5nSvXR98PCW15WW19KyY/2s0+mHcESb07HWQpdU2R+Qu2w9aVP8
p5mV6N+4hIRKPa3gjzF0s0AzIbFoF6khHTya4Bk9dATZ57TvVc9bNFXrhIetsPtwu5qb6UnO++Z/
CWz/cfTgl+v7Xo4Gci41uRDxkzKeksm+tiP14yYO1RI3TGuRubpa+S7XJNabhkt5setAJunEtTb6
4RWMUyGznMosgf3O9TP+88KeiJU3pzPNQpVw8OlJB0jJCaxxa5ZNegBBfw8Bj8FmHs8G/3cWGy8y
4MMnLFVzZYirWCREniwRreOA43clCEztEunsw37X1r94xfQd9J6XDXSNx1Zp0TunMnazWQQ4TeZK
I7EUZ3d1cRf1tuEj4PB6GiBZFObo6ou+785iP6E4kRUN4aTQygK07qgK8aAL8IguXt4Y+0QbMsut
fY5/IYEoGSDqwMwSQEl9/lBKQJAXaGkYfPPFrg0qs1NBKrmEZtgTnG9Mrih0cVHK/HQOk5pMfhmd
2ai7RO5xiUWBi261407+ch9m2pam0L6RvMdsIAEK9+Z5dqGDgy6kK3NqGV7lxa/UUxBC5hCj6nDB
B2+N9Xetk6Wa1drxLDUG5RbEn26qlQ3qy8M6Na5N2KR8EkmedsWulgVRUqWRPjutAJm7Dt62JlVQ
QzF8kRFZsKG+vz3KEv4injhdTWD6uXW6iAwJch+upZmk6A195XWYbFBq1hlJ/ow/NPQ9GwzjpVgt
h7H55it5Oxl2CSv1V9zcDPYMn/gBbSEl0i2AbvSMu+lZXhtKcCtMoKbwZINVqSYAUHVESznroeT2
hcmuyoDUfAbnkFeCM7UsA8BYOeoZ0mkstJDxq8NrV0ZHynUk9jzxXauF9JKThRfBvmWnTTNqIzJn
pb29gvSHk7hXLCznS5uHm37QsK/O83w4+eE7GotiqQ5oqIQE5qu7+RRAuczgREo/UTIjmy84wocX
e9KReZv4jFAKicGd5jlYoKd5RE96B20lnW161P2XQpTa96TuvVwAwFdQYYpaaALEy/hDmwRTp9oj
x2WZlIQb5yn4JPRqE4jSelMtpkVScs4A1qTjFQN1A8I6lDQ+Lg3MiBKeKcLLddt8M/sRrFCLg8ku
rbKj3jp20uHkscs1Ee7yvnMv5AgeghjCBbq+MSHsl4mpwl6NFl/KXRJG/gM6JqIdzyUd7kyuZlTh
5lhzIp41KzcIshZ8/wxMrLDDUGJ6pncfxUQ/dqtEvoTjM6wHrdgxRrnVKMALAb5UPM9PakdklkMM
DawxROVKquTz9YDUJPGqrWliVKbBZZG2NgVb+fBhM2Zh1hfyHmMUxYxS/ZIV8DsYFZ1VUzT3Xo/X
jSt/CQZjA4dSidSzU9XNlPDoWS25Kf4OiDGUQu/ARGbQUIeakV2y/fl5HI9tSyTKNimrDWNnArTA
C7cdo8EIl/kbfLeMRlpRbLtccAekFUO8VQGzcBf61lZ0xfITbtWUEnij4yyeqpXq30hkd/nmHbyd
biJErPeRySTfEteaUrJhm0J3uvMGncRXQOy5SFEWEGzCcP4SxBS29f5Gbb+wF/LmAhVyQOY9Ddqk
lyL+ZpkbHRMAjqp8R6umxgC+6+irt09P26ruw8OKD5C3/45jCsK4ZQnRT9yckP8+tvg9kKZO0GcJ
vWKT/I37M0FYDs5vYSNc31Vo3ENxVLVYVFdFucjCIhDwZy018vRYq4poPsW1K7i0NbMsz3nTBe/a
lr/HdKVFZks4HDmCOUHBu6W50zMhd3cJgI+0CzH2eq5OBPyX9ReHw8GEFLtVufX6E+WLn7R5YeGM
ZTK2d/rjzkjUtRLtRGslaL5F6u0YXFjYAB/gfAaZWadzU6K5VSxNFUCalIa+aD+MXT75Q86pvbyM
MGQ5uUywu6PnkV8830JdMiNErf/m+2VYop4JLbTlPwyXCMsISwqLj3In2FCjp8jQn20pvjrKfjoP
x24Gn5K/iFF+vqDLLQi0q5SRBwWzob9dm/SVG12b9Bk6pTeeMyyHNKishchvOyasWU+eLrV+jyQU
NyPJ33tiEkQoB5UT4msv3eOJhsTHn6Retgppix/czlkJjLn4OjmZsk837nWrFAqn7g27mA5vl3kw
0nx5vuk6O8nIq8uRsy3I579djrbSZFUTZjsv0AknADrMWKUTyFE7gOjl+n1t3Nttc/FkfttlsykY
RiFIp32rgBjFaH0ygLeHR8LYnhop5DKJqUcK0cQ7jL+U6UZgBJGHf6urkgSbzbeycLx62J547Kv1
rv3e8mMvFDr6eHPkdUSuMjAjRoxVnZDWq4o0xuDx47NWioEyl5bTzMSf5ZHDVZRPs7i9m1/5SU9B
7nX9YGFsZHjTWM0ZShP/O6LobyPEG7hM8P/IvI88xMHctYrwrU+LjQW+Jk1JyRxyvKgeJoriword
DXQV7IYhv1lMv87c7WwNpRIw2MdbJYeDZuTocky5Q/cgIQ7CJY3vX9Q/eUJk9UXIrRmF1d7WGyZz
YIcpjM0/uO4rtryF1nUugdvnoPSzsBxtISO4WtPm9WpxDjyRg8iw4BIp+wO4q3pxGcb6l4ML3Lai
GL3grr+iteubkiX2pOtspJeIvRZLVOS8vvn7K9l22VO3GAIS5LxRlFiWS/+AiXTBBrIcplVMB2YY
9y5GoDJGWxiKxJnqNFOQ0jUanNqq9zpim6PRnztCcITj3OiUaFGmGJjeJWOn7BX7xCvNU5JB+Y1H
+x03KqIYXytZgcwv+iovetqTq8afDcOovYN80C/EHu6izJEjU8/mvX9ra4/obMY8Ui+ZPjEZbBZN
TvG4q3vJOg0ZnlnVNxLrGjFgvMIe9engDlDR+YOoq7948Fmtg+zh66PAxheLiyp5LPuz6lH1yqLl
NZITHgvOzpjDDctA5gAcAIpGv/JWcf75FOFkfhiQ+Fy1Rvsren2KWoCffg+f4iZlnf+49J6Wep5I
S2xXDol0goCfw5TAyk3jdAzIVODe4aiF/mXzOJQWF/CfMkIc/8JAOMStu5FqIiKhEGeCgycBm2VQ
w8gfxLaJLnjCVGzI1z5E8bIRF2kIrZP6XOBtI2SpcltKIwupgULLeCPytFtK4tSreStzsgvyvVKr
ktaF8rFFlkAjnqPTqpvPCnNYGhnZBeBzX1smM0VBwjf0rTpmBu/t64MFAMWvqiN8XUrzFq0E4oDG
9uMMlozvLB/bjm1nbNfCnYn8TGQ1NnnhEzruAD+SHju0ktYRGZSjaygHnUlusfat2LWswQat841i
cFOB6F/kg7cgSZ0bnTYoluoMRbhqMT7NnkpPkDqv0+6gzA7gj3V0981rCC9oQg8dvJC9xpeDBISR
pXkxUouLBaKP6v30erGglwnWyIzlGLlqAgPpuFtZdMRUo94IBhSHhIykTowJ9NDjPR+SMRtmsJju
rM5vv91mMDO8G6aC8CYNqBcYKneBC4vDGFU7uhpYVk/OMhF2pIO47QmgqguuGWPZEhmn2drBR6Eu
7oATlo9r0v144hnZFk4McXC4LwsKb5JqoBunSNPUSgUAaFRoiqILnXiRCfSfUM1YtO/iMwffYLfE
f8EUjuKBYt/DJbgEzYwZxwnmafY/uE/ea5ezJthQI3gRJz8tnhVGU27AvLtJ829ge34gk/ju1Uyz
aD/eiyvK5BhgyJr32vHfC2rpN46TmIdZZnm8kjZd3BBF+m+XHOoBgYPKKxRAx0B6zdpL2F2teqmU
Paffm89riuKZBm+3ZcdtTsJ6wEGR5YiWV6U5/vpIDm6ce+SuIU4HLJzx9mOh1/jf1qOYmLfN/Ft9
IimaZhHF/Ises2KeBHRL/1TzTZSsOG6qiefiDATZpmLjZKIvYM0QdaJtMzX7IZVvsvmAOQvD5caX
y9W651fKe/5PyaefvIvp5FpYBtzq10tOFiwyIFa5LUu3m+E4EWw+TgeFvOZWZspb3XiRTRzQo0Vy
KwPQG3YNxVtX6sYOAEvQMjZhzYVcVDcLULxHaLde6SE5aSRuAZwFv6tfcM+sCPD5hmiGMjEc5LBv
N2SBnh5laa9r7C7rqQZimsghqE17xuCvFkLV8b7ehOgoIdMEaywv4Ba75ymNvBV+HGAGQd+3tjxY
HY1b3nSH6LRtGurITxv5GZzdKsJadqaFGoVqwAowkJpqhg2E/6J1i1RuESPXWtFC7UitzmMq8wL2
RK45JGyzBMOILFVvCeP15gis7qhkI5yeJ7Al+LasPuEyFDI1IHQE2y8EkfZgOaoW1tKEgYZXe3X+
BgscW3tyTI6w4/t1swMZLOXnVwj/AWuJlIy79HXVWZ/XGDuOCJ4jAk3H4wtGiwoPQJtJIsz09qer
57qk9ncc1kANXJ++1yebr4yYAD7sp2HnV2TzauxoOl97UMQFAC1dvpAaGJ/uYwpai8Z8FYl8IPdC
lm4BxMcyON6PIvi1CGcREizKaFsyL3SnlDjsUWpbIJ9hlQyMdWF43eCDzN2RyHfI1WMiJ9K/cesP
2RWG7UIFe0iJyhptcdGNlU9a9nkg/BugBeyD5UUPZD5vPRQTU7zx9CD9LJQM7Rdlw4uE8H5i6djj
aXSLjBPqZx8jyWrw0fMQS0V4gdxAdlbyeYsbCn18Sk7LK300dSRS60U4aY9+WewMLby7Z+V7zlYK
DsYwOhXEA8Rq+kfcrhnh5/IQJ6PcmlmR+Dmra+6qpr46vgEbJzijXcwKUzCXAiEW8ZNGdKrt7o1e
NJgGxewK3KqkWMcyfL8RxBWubOk6Z1VRI0ShRCRR5Ieck6PVvlksHI+eKEadQ/MywRSvLpRSOJAs
I3q1Dvfxz5Z/HuNm4vP1WsLL8xVd67pWntNp18p3lgc910EG1wKDU4vGD57B31B1Uili1/8eyhp8
jxr6ecR2xWw+6wa9P44oFTE1d7VGmkdqouKrIkBjacPHRV0q8ARipYl4nIvDt+YDVucGO6cZ9oN+
iCL4OiDTYbH9r9X9atrXPx78Sssh7iY1UD7jy/4Docsd06bdpy7VWu/zpxFaJv7gi2slx8rqgdl0
kl/B6kqCj3FNeeuMYBQzc9vXeXtEdvHf6VGyHDKaJbJyrFytFcMkeB/KH4359B3sskTgFWmaLuYf
nz2WAkxc0Q/FN1rCULkKb1h94O3Twr4mUBb2MNhNjJICMGCXGgMIas+YUsKxxOI9nP8rWj997e4u
WSUYo5NjIH3W/z48XuEt918n0RNdJcPTUK9ETAfGIe9yFgFDLVkUJ6OO1w0y4c20Pxun/4fL15BE
2JS4iwz8Y+My6rW14OsprqNk+P3/5//b5feAA1fZNZEwFkJylrmpE3GvU4CSEgqdcD84vubdJcpy
0I3widfhnq+xB80fivfRriVjnbj/ZYc/XO4TS7c7PlrX1H0pFATauVeRsIZymD0M9h4Iuh1UKNfN
iXDXeOQmPeGJg+mAGxDvS2a9ocrL0FI6p9vpA47LKQUHxYKAVKEP3gtS1fnz8EV6pvYncQbyrB+S
U2kahmZBX0kzR3qQP9BDfEMMSeeVM2o4O3kgJRiPFq5M6iqF0tvjPrG9il2zXseAE9ukQ2/agL6z
roRTUlvK+M8ftmF9/quTx+SOOzwvHkUY0GlvjUN6zkHbBS7pT10afS2Lp+zV1mgp4F6ADpJv3LRP
Z3on6QQ/0oJxjZlmRHCCLW6KQsReFwtgxEDYffIHpmGklWgskz5+vYfj+5dZrnFmqOMToKL5URt8
L29tFofq+rMK8BH/NGm/mWE3pxB1NceAyrMpdTTgAz9xswAT+q9Yhool5HupFRSzo664liBbTSGc
qoF7lC3VcaBHPhz8Wh1Vhlnb/xkcLsfe7xGJFHC6H+PEIZ+aKtXPUehpnMK/NnWl/UTIJI1yJiQT
/d0G/V2uSWoZ+u/Ask323kPKsSr/TCVH7MkqtgfW3+Uf5mtRkGThNiINOJcwACL/qxax7mzvFeI8
dtbf34Zr4p8rSkceBSsJTyLyUD7GLAi9Z1By2ILNS6GBZQwXdQYEcNLEwKoESrugEQPIozDOFNyq
VBn81Qakx+G3hcDtt3RlFOQ6GGAt7FuwWeLfzU1YZfmXjqbwn2SL+kyXHLOssjhtyvz2OTivDF/V
wF3FjRPuYxIeA1gou4//ir5M10NCfJRphGFuGMErILA279DKDqKS1Ld11S7UzonlLqDVA1ZN4ta7
wzxUwHb3bq/lR2/ZkOtdcvdQFthVoDE/0piSSjk8madhPBuXn4KkIodPycHM4I8oTI2xuDouR3hr
Gk54TE1cEfwU01A6RC5wDXGkx15WAfrGe2BOgOXqn0WrjWmuhqPMbxf1l+P8elPAFhzoswFHNT2i
FIfTQVVD9K108+JB0HoblbsNMcjofBUMuSUn1QEHLPPBNlX/u49Hv3RJvqRXT6eSQQ/6NM7shI73
MRaf+2UEjqsH5Oh/xd1Q7Xs34Lge1+IWNJNLzL+Hy9Pf6EqKT7HhPT31sUz1ABgON4Ryx2VIxL5A
A0DKbnzJg4gFoKSvYlyMo1j6nv3Ihp/U5uXOKQsryiDdG2kVphJ9gIH4pGorkODvtXUR2p4/o+rw
RZzp4oAi8Ii8xsYdFxU8vYKMRKsEDvt8Cn6mvHvdo/uDqOx0C+6n5YN9qHipFotACMfT9HV+Q29q
vX4vN75JmLc1BA181+y8MalGYYVU1JAkF+QdkaYtlyc9MUvJrKFzLgIIUffxrFP5+++Hs+bm1NWh
enmj5gaPothnYmA3jdWUwU2mAqO91PXQEFdPi2CyfNnBmunazXePbvODbETupsFSMQv/mrF3ssw/
BMV8Yg0Frx3huXiGS7vIUQsacN4EWFA92Zpttvg+QMrX/NZdBKwnjAzdZICNhuJYs/0zk1J1qO2F
M3GDgkQzivj2MpXdz2+EA8Th/N1InZQGKkwyK++KoItKQ+Qu08s5EirXVdHiiMYd//SGrxoVk9Hl
TSih2vl63jrx4VmBkTOQyRlK9K83rpMcLvW1YqQuQoqaCO0oDLRba0LBWJ5nKazxnUMj9j9S8yZ1
tEpdRqgt1v1x/bx+bwUqX/d0tQSgftc0PY2KqmEeQdI5jFm91JSD+FNbeZpz9hf07LmKkxWbFYmI
D+qzJ07P3w1sK3GdKbapGGwk8s81HqJ0L6T+EKGPGEAqMGJD9gzn3Z1MVCWubcfqjF2+04yhslAN
ML+I30enPz69gjweSNbnEqFwnhzl9esS7BevX/X/+uPTEDbZJiaFgNL4erylZj7+JWlzPxAFq9b+
CFJhV4NArfmBuC4UDt7sZji1L9MZAvPd4tMUMauZ0CRRElBT9nDebfmze+ki60FFdtCZ0FTBTbkB
VZohJpnV+u6n6cRcQtWaOU2wo7ahUJySBe0wrUFFu2ORfhB9nb+2U/mpNH5L8holwC4cUCqjPQ3s
7Li1uX9XzFA0ZXhMN1fxzy9qjQwj8cheGum9acUNhPt9r5pLeqKbG49ASDew6znDmu+2bbxfki4+
d7aaJMLNH6W8BGb4WejQyW37qEJB0/a7L04DnhQU+1c2RDtnGfmM6FfBTgl3Kf10tN0ir8JeHUJC
zjq/nWzliXIn+Uxf7VxeuL8BQItRBOXZp6A/j/FrnjR4MZo/EodIk7MttZL4Jpp7BthuKHX/JSc8
Yswsv3HyPcjd719qLzMTbA3o+HJ5ziKUIg6TRVHCc//gDvu7WFWad7mywxYu8256a7eJRUXBlAN9
NG+st2f22f8a7SswyeJ9t2hTb8iC1maxeQ2PFycuG13DUJQiPqirMoWGpQU69G+E/+SH48Lrk+qV
/noWVTBiRzY8caStvWukpCmNwR9PvEafkc6+xzEZmQXRw3xeMHI6TcbLyIX5vQ81l+vHB449NeqG
jK4+vRafAuEb5cv45aDaLDADQfAjTINQPn5hsxRy0gYusXZy6KRcUE9+wcaUtSETRNVUjDHsSnF2
iJiBYI6EcLR8tG52eI6OcY/+IuMs+X6zTQqIH/pn0LC1Nd941kTM4xAIEJbKQcJKpsmC3BwhOQhD
ZCHiVwL2h/6VgehAhuSoAva+ctDafypekWGIb4/nfTgUUE8Bz/i6GlOlRVog5U/dPFgHe/lOaBUg
Bt3731/PxMKOWTKyj6OS7FhVSoNfdBgVnG3F30v7KRvbziPxG/eqMptny7r8QrPly//WclcuiFea
bU9lxKEZuBrwgO8mLbLNS3cw/bml9gTsGg6aXz0e0Ywua5JSQSwca9HcxwQlPRma3/NPSL4nXivY
vwYPRTXepAX6MTsaDpxSWFWm8NUyxQSB9o18i8WnM0wdAr9uJS28keLxgwk1dyX1cQ/cj3PFKk0k
z8pm5v+jCxJ6aKf6UpNKZnNb0U194tP/B9KUQ0HQJdjXoiAYdAeUCq0IvUe9k/Jq0cjG4vlRBHHL
H3LM+0PNrLgXFEw9FnSydTfmEszn+/ID3KFum/naJz+4zF90yQxT1c7Jvi3JMVGzsJbJxY6fjWQb
ySnGVBYf9a2pD2VNyZc/zlLOCgbOMlRfnAgzCVoTy6SyMkUJDPwreFAJdp02xqVRm9WBPBAATW8V
UgiNSR7BzDNUhQGKVgH4G59oj5TM9z0er/jKp5ZqHeLaorH3L4Z+WBhs4/i9RMibhyjIFZx30wfe
wTKzffUGNAFb8NpkvbXwN8BoKmaVFIxYCfkPZgKGQ+mTpy+saEn3n9WtokFv5w4UHn9t0e5L9MId
8oOnLbDLBz27FVG/wk6GZZxxTlTxf0WQWEi9CSj8XlXzF6oWT0p2YzcrmRkT1HTfV1jN4FX6TKGi
H1h0BvpOchqioWuU4nFDZ1riTzMzU/ZC1rdBj1ZJ6GGH+vjFK/ew3gFzITkO+P2JPYuY6djUod8w
xfn7kIcPwib3YsZ/mySYGbNDkvJKFpClt2RQINeM9odi17sP+3nmNzGHMrHYTYWOThdRcx8LbuqJ
kxo7k/2gL5o10AkOTk3hlwCvQMcp3p3BW7EEKv4wPcZ0WDafPFjZ3+dXjiR/MfnHEF4Hlprh31cP
JHcnKRkAxUnz5Ho6YACAbnQuHE2s2/bHgbsKNDVEPxK2u0zU/c/DMP5GAPiky5owp9HgZ7Wf0qC2
y5DHg4R+D+Wj7lbAC93YRHfUDOA4zLeJy+UcSQi4JFJCTO60w/tFs2rLkeeh8vAQ1cJH2e02YJsH
qXMOmB5nKDRPTzFoAuxyGgPI3UCqnMvjcOv8qH++BFUzAMo5F4/PHxwiFnuLk9/I1wTMhybqqSUW
ZnnXb6JcVSeIx20AJPT0NzDkOzpnfX5tgJUedcRtDtDpPALSoTCy030srhWgMrH2eilg5sed7/Uo
rkCoVTFIhoj3jhCf1pZN002/46gLc/8mdYC0hJVHiPaUQ+abepVc1EZN3FUP9tXbjUUTgdk/1Iqy
6fT1KwSt1VDhfA9yLXOW8l6V1n7iWn3JERazsd78jXF/MeF5iRdipDTZZE2JdtCuCP2Yo/Ycop90
Hi3/RyVsvCgrjfc7zdWVrQBBC30o2Rf0Y1CECWFWul7TONoDke2yit4LErRZhtd+UAswXCF3fr3y
A4MmfdGCjyuPyRw44Y2Ip7bjPGuDLw5iccMzKKzortiRzBPMLYsyKFSgK+2U36xspPz9YkrB0thN
gWLkF/5XPjZ7/6descANq2VcKsEXSp/J0FJOLwVAlxmjlcNLocgclhh35ch5sFClNxsncIs/KIEv
EX/831OggYPQbfMKum9GDVMV0gKQfR/SKSNZh8ITwlkmVxGN0av4WpamBb14JqANFOU6uWFAh4cC
shOoWEPBlxnxqU5YbqM1uB7Vb7cfiomeuQ+5WUkCj40tGBWTcWcqv3foHAxGWC2+9eV2K8C+e6NC
+TbpqgMM9kIgKPyplPweUaP/zh88g8W4h8BvMpotYJzm4JbmUE3u9gxrE3DDq3Z0KRXy+R5Gl9Ch
cvHFT2Inmm9DgJmuc+EKlbKNTa7O3+HN28KmsRCuqB9W0GyfUZ3B1BVZIz6hLnoYpWB5yUG0KGhy
d+9vsQzREV2SzJbCF2LCPRq5LyUIYU2LlSlg99eYmLHHaqWBXZA5ZvPOtGocbWZoIEMQXARhrm4Z
MhAIub7HKF5Quz7/IlxjD5sXhM9UyQoTWgJl8jmBBSsYHmwVlWR55I5YyL3Yzgyvnp/SYTWZNJ/y
+TqUsGXJI5fOerNSGf/+oEikw7ClJQnq/qqEvGmuQ1Q9BUt46sHUrzqCEdIKBzzU6jJMj1dJS29Q
8De1tbZYrs/mQxnmtJ7lzypo1T6pqj9KWVOz8CqzkpSg7G1RQ2iGN/O7NeL1K9E0BUQkLzOo0v18
ImeIwk8iToqiN49GssgKx8rL8LZr/QLTiVvYHiOz20QpgFBkuusbjWbFGLyT7sa2CIHdbO8/4uYM
hr+Pw3+IlJWMrgBasZqUwRKpuZW7qfUVjfQYswWu3l2Vz28MpfABg9Oay92W7GjA+Phe8brYmYc7
qVMOsWrld5aFizHxpKT6YASRhCpKGBnjv/hEgpwu5t1sKUi1nxR8T1dVxGhvKqfisf9WBUgFGu5H
gzJKj2NB9bIvFTvZVcn813VW5RplKLibkSv2RkW/a1VwwAl5Lxxutw8Kkd3xdCjOihwyviG2HuaN
ZhRDv1/RXlJS0JNPLwVGK/1BD1Ay4bLCZRwDvODRfQwDMJ9qpY74VfRl2lmcyQdNnIzcKRw0jVZ3
ZTRwblP5FaSFoUVe6THjJ7NDYLTBhDE+d9QwkHktzrLLHFleOGuc9eX0dukSpGu7ND6AM/1MVheN
rQbscQbGt+jnbuGpBG5UFHgz88Y44jBHLJByuDu1cJKjmirom0b0wwmr9wfjmbyDPMCmdwg6mndz
6eDcbyMFTiofwp8QQVk6VV3nXXpBbES2cxZgIdXnag0eQvwdekKnyWFseRF1yc9GkihJWDvZi7/O
Fn+eo+fl4mfT9X7sXxn+zZqLYpD1JYRGOfQV5jJp3WdWHhi1NP/U+V7EkRr8JXX4HIXb7LYSlELU
QFaEh9WPhlniU4dbkQeS4w1mKo6z3NrRxXddNIGoKMWu6nWJwYamwqfUbnT/Eh/0DAzF/gdQQPhX
k76baby62FMTcvCfHfBWb9dU7tuKXtFc5WlX9GQIVZbD+zDETjX8pLj5r6IJnYpotEQX2NgZ9kAC
wbhiz6mNqRtUrAiVKCwFoHgsmYmRjKETiT4uDvt/srISMrxs5JMe88c+0KpwShPTogk7OmY+UnEz
ufnyQnD3/jOiH1e9Z9CCkUaU3tCzBGAREQbWA2I8D8Z8M/5IuzMVrPznHqRvmSKeIcKEVdAhHF7J
IMEJNnzbOTCOKdNHuUhWAZrk9j1FjtNwkON3UAHnvC8FmnkyIvwZJr/Ef0b4cDRwUmo6gmnICCD0
J9G+eIwa99U49I4PaikNfhtWacbLdnvUJ+X3mkkku7u/aFYHXw/QJBUnxdDkks2MSMqX31ryd6Rz
O2U0AZ5nPye7QlsOOtPbhUHjY34PmpEFwPv/s5Fxlbtt++wvfzDPc1+WQNWRLYApRbl0CooZFsLi
YYuLJ+QftwCk37Ba0G9XRsflrQSm6Arg9D93EmduaNUGSI+7AVlvfVul6Qt4dmZsVbThw0YnTeg9
cx0lZYF4RdQXzyDeDCOgqz3esVcSE3ki1n83hWz8TafWk8/dBmk+JGdXnVUgyi+6nLqjPfIW/epD
swsF6VJjxFpu5XnbOEmoUjfZ5xZ3pu1XRMA4Ss738awfXpkfjYaWk9ZInfSURq9UXCdzbeMc5GYy
rpeQma/HofZFlzCJWnPca1Zdh6eGbdNxL+JGfyKi/tU5ot7DzEXMaTY86HDeiowz7NCsTkSqaU+t
JpRvxhB3NQ7qIACi6eOrNNcJZIj2a8I+prGV12jUmHk18Sx3cWhLTFnEh9atMIHyTQyh9awYPwIq
K4VqOzAhKg0rzjF0fnLpUhD0TTPgsGxf5lYJqSvecQg+Noi5x5BWaRzZtBbhLCfniwnz7N/emLW0
T4aMx1MSVyXSeviHHjzyoLzW0u4qKuZH8F6ZHhRp7yh3t3FWlhd+elD+AlIg7w52vnpej8+xKPTu
LCKWtc/Cvp9XJ/21Ry95GHjsu1zyKp+cfiRnkS3U0aKPesYnxZ6tykyzb0F8gUYaaNJgAm8yuRai
Cx7YErHDvdrxl3nsVzhWyWe2J7MaRWVurWPwtkgdJDyPZFYUMR0fvfPhEFKIBgDF/eFji9T+q1UL
LuubMQ1MJEGlwmp0a5gfPrsxJrrmvSxK4wRYBTx6317mQn/dbcre/zFbQoEBFw20MPUegbTlRnwu
QbHG4TwQ0lT3cUR/HuW7CG+88PFc4FIPGKcn3rgnJqOjhDGnhHM8TIUneLsMlpD+UenGYqzUn8l/
7X3Qg4MNlsTl2BfVPl1kOtCk9Bq0Dc0WyU+EB+1ScSLBVCtKzhyx9Jn7+bQstg1iXsmdLGv7RFvp
NBfp94Zch3jkZkEitN/XiOzuDd4kRl64dl126ZaFKkjhijAo5JjcKJp1csmb8fln6KFXbM6s1qAf
kOEmQ+HO8jC1WNCbzwvJ17/we86obd69sVo6bQm6C6XY6f50rZjQFQbv3RArlDxP5knEyd1Od+3q
2FguA8iahHFYIlToUjx7va2UnnKlVKOia1o2fJEMiuBr6k5pBB8kQBfEf6zyi7ou+MKAqhzGzCzB
iRXq7E3h06+qJHGGSIQIJjDwNvnmt+Bzi493tsqn9BYPbUdjaSO4HaqX3ql1y988CsFRUiK73Dyz
VClNrhC101dklC+rmkZ6Felrqr2ogsi3BSNY7td7t3d40DWNaIJ5Jo+8zxwBHGfBIg1R/strDQgd
sAONhBlzC0WO6BJ99OZW5LIXmxC4/ZtGzVqlWEdAwGFjIOqFQDl49LjwBDUZasTs4RXn7sJH2osw
wT+TAzjr40oQRsby+ItoiLUnX8OtfPuAoAk5dWr4qi47/oRcEtEnXsxr2AaWLpF0nwBX2dFR7KXF
LuSa/mpVg3XOSwHeNfexDHg4AHqskzOkSuKoKVjCUyDFnCgpJjC0yI1KthNLEyUW2g/Eie3OwoHC
+jUT2tso93mQsdOc1TYwjksFxoEVRRFoLOWoimCCf/lxBD0E7pURulQAporZKkc6M32F3TMXjyph
DA63EDfPlcZwrCCLGNQ5GTq8EwRo6HA5H5jJz0N52C+9YRmvZJjLgXF7J+WlzYAhYcNF5AXryfb7
J4Xe4UmkzmxYTCgwAJmozFf1TzM0YZRQ1hTcrDMP2I4uQdux2kqmAhUr8Pj3OrheV1YHowpoOjuR
0u9JD7pN7CeabI+ScD9yysfDFyG1M6gnmpf0Whwa1SfzkOvSrNd+WPOGtkD62MxUem6poNfAPWbT
rznJi8XnQjn4etGqfSBetElV4D4Ary2jnS+X27PKiEl+T/98xWCF1hTuQM6iqO/xCCn+MbkjFy2h
x791Vnkg5afOCZ6BoM4bdio+iqxc+ZPjf3osO2IzznwuHme0SXyJdDHryBjg669lL8/SjdcHMT4X
qBZWKNHiKc4c6gG+/R8lWM1xh399V+dZnRaLtACIN3VvRRa32eHW0NooWY12RXUGye+uLnFskPE3
Wdaw9yIg6gtXTB2F3GHaIhHEtxY2bKirdn2q+FL4FYdXCqIQvTdN25UStLPtsMNJRVofzzCZf1CS
AYaAghdlfTveBzJPwfSn6JWzKRr00w3EPsif52PtSVHBNs14gWqBT3ZdK2ZQa/PLz/I1x6ZlMHwp
bwFgBeZNIZ4qDYbxxbFTeBm9xigY1TZI2mLFtgAviS/JTHvIQkRh4EHnhjGgu+xo5BLI+GAXvXzL
T0WHcCJjGuOqaZjsJrReSGCgKcQeHH1Rr+xnOiZXvzefyg+c80wMzKQ67a6w0BJN+N3uXknYA8Vw
5xIU7SdL2wkLlYGnmO0DIsZVWk7nH1VpD0eImGv55f+6Y8mp0H/EtibQPJvt27+4R6m6bnaXVdFu
smxe4jB8ZgJcsVcC5+rGY+2t+vbTYp/wtirQ0cYSAVMmZPqoOisXjTw5qaTnbeMm0bLebmPRA4rt
btgKdamdGsIIoi3aZ9kRaDjzQC8Xy1LEA7oijDItpk1i98Dvr5RupverkdRC9KI3iLvVRGaeqUIT
wfrjFRAeBvjOo3PIO6P/kmulfOFbUWRIfy5l1oEcHvqLLwn0BGqv2e1JjOG9tEwtRx0D1OIXVtzm
zPkDXjclTYLkNpbN/el/E0wzZE4gsEYgKQDVUPQworSZDq5/vb3IbtxRgPnE4N4355+2wi8cBxVS
I9SY0zLX/KD2OZB4FCX5VemFIiMwyNNPQlECGRAtzzUuo33WYsCDdAL2hg8+fTto+fyKbynS1g9z
mrmWTI8gzH4bgNirvJ8Kk860/P7XLFM5YwGoGQgdHPtRPU+e+tR8MxFbxvKFtNL0nlboUboyI9N3
kMikYz1BT6cwRE8Y4fXpq9NLlGTO4MjxA2vOvRiB+N2kvnCOIatGfUVsnMOEmCP5+jHij1tbkJMn
w17fpF53OJ+d4HSNibjTeYj2Wwe7G8RGjnD1sgTJiHBSlGqhVoiOURZ/0z50XCQ7+01bXzj5T7Go
lhuWSRQagSHzKLsSvko9jHgfCSzC7L6wq14xaKpbeoiPIa0tQXUuSNpZdNbjGJjaO1LG3pBRPEad
yBfw4sIYi0PYWdM4bFKynt4TXR3dXA2ZYvXp8OC7qrL/gpqM5Mg765f7Nv5KcLxZgf7gDU4VcHff
tjmUUw5NuRmfH1MTtOqt1dXBYy3IgVSGDmDUHATDN7sm2HPGQUTJCIfTnbl43qmpP7hbIEW0enal
tVwSpDzyGeF9SxJUMedo2I9R0N0X1TXsg99L8D5zHjmDPNOEHz9xuX4uXz+oqSAg8D6TxTXmv4Y5
ItP6EdETz+F9Ib+Z56F6hNBzYCosXb6paniFoUdeIdG67CGigsAJ+KsEbzltOsQVOx9OvXn7MPq3
BUejQwBSmcRpM3EDSn3e5EYAen8MBsAIjVetLm2G4OE4/d1QjcDLbq5jAHCx7Wsuw4ebxwoayZzD
1wa9CLCfBmdF9IHODGgKq1qlyzLldRsI+wSOVSa7ODRdJxcVyGQt/AF6zln1NPUhmxrmiIqcuMo8
xDhHNibWlwHq405EvMs61E7BXL0xl/5HJlBn+7R9bOAahuwOXRb36i+ppMAJZa8X6VjOjDgHeFtC
DZo+fWdeRz+020NPX87ebKIdOwU2nOc6UALdyKIFlvZk+Vn1c47gC6hjtHYa8u0FuuhNuM1FL2VJ
go8jE1CSMpOn23EGL6+PSYD7SGg/H0ZhrRDoXumm+4swr+6WdlJkVJ7CpAThW+7Vq9HvwfsehlNn
e76VwEEoVlQV+hT3ozwC3i1kadWmTM91kONwYRHYI7O4iMlG5wyY1QZlZ7/tYP+riwgB6JAf2YvM
ZJhrHWnu8SQNFId4CJp5JZzN8XZutLG39TMeVzmc8ud8XPke1zIhAYJIkYbuxo/6I0cmT/SqpOPw
G8bKKjLckKG3FP10ays34gLZRMel591ZOKp2yKJRPJeDVEPN0vsFPqgAtrQPJUMp3JThlklF8xyo
9p3L3IrwK28mQViRmGpRIczkXOebeP1pHMDzDAbP1bWv5bXNkZHK1hFF/M+o7JzZc5S3PGFFZ0Tm
+74t7F6qiuQ7oBSmrVLIX0tAQAGqVNWX4OqAoUzmlr2YOAzuHrs4GTB9diFmTkbXifct7Jr8P3GR
srmQOWYsy4QSpulBq1hfDd8i98XNdUaCOTqQ75dgSP6PP7DMkh+TlEolnDp51V/KGUdzn/F6dBQ6
HaMdLviayN/H60p8iqCtq2B23/WqdViLutLw/XjOsl7C8RtodxdZdLFcG4s0sJRlerZz+iFSnorA
dWmjYGfflpDHA6Z7dA2wjxBtgpM6sHJbymkKxT766mo4HhJrL/G6brBzQmY5JqmYXwXrTnG9M9ev
4CqUdrfxfTnohJ1AvPxZ2Hpxobpv+6fsb3+KXDKbm8EMh0RueHZjcF28hv2sC8In/eaDfP79Cbf0
8P8E4KOte5qbTaIp6hVFh9j0uV5/QYUpql3nYDW9HndTZhyfU2zu9hnP4tMkJnEFWDCyEVzSO7XF
5zcQ+J2p5A8PT8d9w34brLEp+/uDO0yDIBdAMx8nWQ7JpA5WFTuwiUQpVgjgMYq/BKhB0zSsqf6u
u5CL/3UmuNjSkLmr6iIdy1BXDVXzTQpLjXOmpj97m2bLuEuSQmNkbfFkQUmKabPMmwY0Y+vwrAfn
HYjZqXmCj+rzls+ikesxlXl+zElI52im48T4GiNGY77Vz3KUfCs7MkfYUEYvJtZ77khd3YJXsbwL
8XrtMCzuZUdN5gW9VczGCp7BxGPsQjFZ/J+AjnCkiAUZFsE7QTZLTiDxZef7UH9wLNNihzZu1fsC
PjclQZ3qvQnT2f4GEQDdATuYTAPSMWtqi9zvpuqoRLWLrmB9nUUdI5Garj5nTus4QSJydTe6KZXj
1ttxSAzggYoSIml/xD62yx/fIjzc3W2FEFj3xN2K0vkQR3D6pv/Ew5T9vjEbWz5zDfhMgGNubD3z
D82bsQTCblfpyHiBR3JhtjbOR7vA5tNfAymqX2YaafisznpyewEzsKXWfqium8/SH6ztvsvawARj
ZHEyvT/hjwsJtdVufQeNiLuCPsuR2F+SMb+pBMLvYq1TKaQdibhL0oaCtZUm/sw4Ae83rMbOGXdn
q2cmuc9SKK2nyGETua6YZ7S540tiF4r87g43z/VqHC6oF811JlsQfOCjAy1FMlgaH3XIoujXhQpG
9wOLF2qlvlxBRfSPI0YFBXac5MA8vlWa4bpftwnPjy/xGNC0gHTx3m0fZOqbNkDiAdmKaL2BbvxD
V3e6DcZX4iVj/4ArwsES5l0YyRzRWRN4V24kuR+XkgZROzvamZZY5eCcGni+RATcYodbWUYhVr8G
+vwOB0WZEROUi9vEHs+XojsE/LGw2qsuH7phtsvkPRSYk0bOBO4QZ1kqe6YWdRg/hET81iMPa5cr
eDOG8r8T+9tiArQfCuAHedv5TKp3TzyKfvoZz/iGv8tUI4T2U/oaSLBRltvCIL7aN9i3Qlxk4WwU
gPLEAg2/WVjIxYGkAM/M6V7ntscM47oXlJGPr0ZVQDzTtqhMAKSHCRf7eDggYPIFlXZiUw/UlRw+
ttBVUDkDDoEx7dfIIU7Q+UDC+BEEJcVv5W7nxGlRMnoafcOuaK/a4aPutJ8DWW/RcpIxMYlPwD4n
L+4VREVMiKNSw3NRhpGocIhjFJ74Ouh+s5pXIXOjS0Sq03ep5x+rVoq6oWsAMU2VNAdyina6Rv3v
dVnAWqO5b81qR7F1lEd52JiC+JNSKIX4lANXX0CySQWop0c9FcQUuZfB0vYCShRIFhbWY7VVGVJr
Z+6a+ezODAJO4cXfGgX5EZQ8pchw53WnDHzcmHS7ug+JyQQxsbDgXELEMK+Z6zkQ6puXAtSoncns
tBoK4R3W7eegMYmz5ABr/6OqkEZ15PoWDwOhoElILVrKg3UjcfhR3rVQKgMFfn/Bq30yxyRgMSrG
FIP24Xb0p13d20i+P8ADCRqnI5l+xAV+0fzHi1puvlt2Eg6QMyHMTaD3QFveIhCGMaGLTWDO04oV
pQ+U4ia1x29ViiA4WVs4bw/hnzIRtzhRMti7cwTRfhvccgsmrlpYPG23p2EgW3zulUWz9UUtmkgS
sVhptVu52K7HtjkmqhwVaLSQsqd1uwzBXjsq7L67Qh9vkgEPCNMT2lxnAx9U3xAD0EzCMAJ/zYeV
5E6NZE+WoM53Gy4+c6wGE7OV0VV99QUC/eWb1DIo5v0r+8g0h6U037nAKIWFPirLt5vFPuan66dg
JPEYm75A84MZdoTrJhkjbjRnbNZh6i7u7Hm1ItCVVxZA+ksS7bPwXNIvyzyGpGCFj9Ncj3yfjRhy
C3vwdemTQeoSK+MT85TEQULugeglUCB+SyssjmvPUZvoxq6fKKUFxlYMhqH2T4YjNWIqK+7pxiOu
LJjZ/9++7rUhsL2AbSGHhRibwtlBc1NBBtUBjEDO74YP8Xd0ZZFpbQw2e4n7Af5YkLpUoHJItgKa
nRdlJk5iEY87PdTlk6ViY9VuxN+SaVEjzVx25iYL1uZT1WGr9CB9jGuGbYranIjd/u0MSjWXheqJ
aNgduP8H17SmibjyMMLm71fsqEp9ArZvLaF6yp6sONKWC0kbB7+HtM59VHR4bB7WSkFLArz2lntg
rXPcsS9kON/iGNDuL2E+PA8dDdEgDl2f1O6K4gUyUyytZV62h6TLfPPz6ciD9JbSIXVzQu6m0Uwo
lIZvt49GDY+LbrqAuWtGkn/6IiSqJYL9Eo5IKt5g53JZGpXBaK42WjAygFfsBeLJii4bW1RHNTUg
Aq4KHC+9hGf8udK+6KMlklDH4N5lV+8yjoeaG2FIcLmczIHOxtT2wxDyrakaUZmlg/mCUd+d85Gd
EqHBN+AET2YvkUACBi8W+XWoiJl53zMXZqJaAUqOilqMZRAPO/n06I44LYpeybE2Evp0cZzV8Gol
+tN/BD43XS9csg1nnEh7+AhIDLkfYPkYXnACgcYIQlpD6Ji3deJmmJp65fR523ds8Q0aoMVcM/8J
q8/WNnYqdPfRa4L83S4wNq8DTEISxOQog8uzhLRdnTc+qMpE8Qz1KlN3LHUbCMCQgL7rTM/2Q5bY
An1Uj/zuOFc7y6ANI2CvySceLVUGn1Z1LtfVQO5nCmmWRwxsWxzhUiOA4aB6xctAxDDjnZ7H3CRi
Di5pmegGwBUPa+q8+aMl6zY8o5iJ8i23LL4H21s9UFCWoBEbKY0RlCCrGOg0oM7u1A0UMdAttz5w
n8mtWyAX9XMbXPRfHJVi3Oz+xqdoEoFj0g+0cweXq5+YrC6DN7tPJFWqmD34zf/xAyApsUJsPV4a
tb+jReH3AXNYKSF995dmohFyEeqomXYoT6cdmeD6ePmsEoK3Rp2LWLEG6YMDU9MqKY7KOtaCxHNp
I7S9mUu1jSB1w96TTbpOZOe/N0GUrOU8DPYjPB/UcHM65IG+Z/geM7VHuNWmH/5mEno0kTRLGG39
ToDASlBkhEPLhGzuj1aIN5ebi/vxwBUBXg3DIPs5Y0Gsxr4gZKVlSTdQjUGdWQDd+p2apGZXiuLk
al9KQIOzmgmpQ9J0WoPwDKYWTPq/WO54UFBfTrcAr4FFc7dPQqNn7mCNYnC3+VO5+tocDaoxggNg
PSDH73rIIaGliZUS5a+Obhfh1Jfk8j6LQvCK4CGtnz2yU6OLuKYW0K5Qe+XNI4vH02dFbgdgYwnn
7NqxFFTirrzGyIxV5HFDGy6j4p2ZRrBrr9xAAOimJ6ueeWbxSRZ4umDz+l5zZrtUzSgX+GUuz2Tx
Z2AAC/SH+83yfe59s4glbFZ2OEF63WyhMtkY4q23M/O65TptN5zfcgH614AV4pTBSWo5JE61g47U
O68ROGQpN0F7Oky1doYFwo5Uwz4t3qNI573wOCkWxgwxOt98GsatdzEv6VFZ+4hWGj0BhkNGaXx0
evMfVxXUOd332AkmktayVBYgaHg8SL05i1BVWAx235tRZ7S0VcQ7PDM2THN25fL0KxPzDxPwOYu9
rLcwezN4D30ta1TEvShJwM0HkgMDZFfHmmKflF5eg0NI+F+YnBE5DvVkuEu+PrWAu8VnEnzlgr0g
8TtOc+ydrvTfC2jAMpugIGXupNUhj+Nuf2+25pu9jPaMImU11aZxs63yiRdYEMsvsWd7C4v7wQmL
5TLJGxFnd/BIxHYHTWsT1PtR0FrPSlhkY7nnWrDMqBDeS/fgp0U7u0BJINTqZgxOABEWyyiNBjdx
sS2Bmkj1Dyrugo8m1BAYwmFpHT902rzw+/tUOjM54BUwsY7N/YMlZFmg808dD2TixJmcGsifSdSE
gpQPyJ1tT5kKJrcbSiQOb2fAnzchgunGpAoz1nB3BAggHmivl5OWDRwg/BdEoxNLRMFgvtqE5glg
LEe4MWic7mXrmNtHEZjnJGOoSJlJmXqcg8qf1UfeyylFj4oM4Qfmvlg4s/eoC3at3gu+erzSMrMH
3CuUVe0jgqr3Qj3juPXiuB/BYWt15jQmfoJwLrYtP5ZUgWC0Jpm+SgPIcm1gIBW3qlkAIq4aJo0m
vyBAcuJoht0Z/FOCsOOuKoWdCjic7zkdyAu/0uxps549io0hVYjIL5DQUFDVaywFzCqc0cJqlUdY
wSbkWWHoHFFCjm+qhK/iwfmkuxSwXu+Yt5uCoGJmxwiffIQZWLKzDFm5SiEgyozgwNk2N4vHrCb5
oJkPIrvqvaPwqgqEe6gsk43F9joZ/lukKKAGYwu2UtPCFcVnLB/QSmG9Y3LZ3gd3iJ42PhYiK6Fb
06rdkSXlSnNjpumUHiGMp1L+zImOX62HLcWsrQxuJnGr8JH7qsMxnYVwgKuqFxR5o3yfnFaBDhAQ
B4N4TDhFun9KW6MbklBcP+cvguthkJ/FyNI/ezFMonQwkiX28UjomfixOHKUoMeK8Lv1I6bN8NVX
aBxaiA9+gCUnWIDDGawZ82zp5jokB6Jmn6mAwN3FoLOD+c0tf7WEU3PjqQO/bKT1ioIkbhtOnVjt
jkJLrPPxZushtqzwB2dhHjj+wUQPbFGJBhoFfYadH6weuGVtH0rz2Li08TF5UJE495n3Q+KmOnlN
yqzUfOSDBH0ftoMn9vtFrRgwjW4HO/a7H5sBxLZkuoGQ5hLF2Cw+MBHGxKeCxht3FPud3BGjk3HZ
0bPwifxHgSgwExA34ZDySvkwZvAN4fy5AHxAUvAfo7Vw0RSXOvsu2cgV4PTCR2nXlOrV3cY/ExYx
8yikZAiOs662TWNDNXLuAgFciIhuyRnYQjpmm1og136HMq+tABg221+HOmBOLoHw9fKpReDp7/9p
IhPLLxku0ZpmpJjc3K1A4Fdx8OFvug3ARJgD2SZTJjZhrQ0lgx2O807m9CJaFiVlfZw9wer0pT2W
ZRebUW/uRGe6AulMFuCuHiBBukwxz7d/L6tm4nhkyJG5ynAJbGSB1cEvhPSrQosbnm0xnG0ehfM+
JIonNKf8678AWO8kGt8Jbet5aiXbdO94LgglHCh8UTMO0paTJfien97anDJMWHmz0FjGVad0hBAR
NRjt33j9UKnhRuXL6lclkgRMMbiajWIjj8Lgb7abEGBztUIY+nUg6kcO8YZTaiNo1FehL0TLLLhA
Air1Fgpt+bLYJzW0TXerQtE2uq45gnE3ykJEQqvuvxNzw3iV7u8P+bqmUyxha7Q0R6ASAjap6GTN
WqwPzYnWJ6R2CnJ3HAMUxlA+TRBIMKAfsxd71cDuT3sR+G/rnliR+s2LyDG0hQTO8UmA4WMW4Rwc
znYv78ymDuDOA+MS75fMF6rF+PsYtptN6p3TINQ3z20RmNZ8pmRYHzN5FUaClS3DCyHSL9fLfsQN
tAXfLOWojAEz3tTjmZJynqstYajYn3S9aMIW92Xrcw/Rhu4Cr2zr+yFBYttS2ru5BBxZfbZY9SmW
BM4rehkldvkCEWVQq22geKdGcANG6vZnTUAfNXmgUTRexbpcjr97ZPq6SLhiryFmXVJt1ZBLDs+T
g1ufLKyCzJsNYvoPTm0F+ldFrGmmCYFUbWH1ryjaO1+sC8mlrd7Ip0mqI18LwcZ5AGMB2OEAqoGC
ZHB3T3lYjC7L/i+tsHicgbU85mEpfwStF2eXzEnnVzs0VyPUHzSye3041ouvDk2+ntemG5YhRLbx
COh2u/vF6pBhy1e9FJpsovQb4+ZG8hDSCOnNgvHlXHxmQat46z9iS2Bq+KMP2ZkGeVWwZCCD2207
zqXwEgcitMRXfM/FejRw1l+r9coCOwEsLXfc7kTcN55DuPsS3Cq8k5/jW9e30sqz7R+5+hammwW5
D4shSoBtnDq6maFp7LAWGIUEDg/73sHK8QyVSnKGcK46LlIJKPEhGQNYdld/08AzYRkrVeTjRsji
Jg3c+/tYgYFBqPqyiJHkk+RG5cQ35jAjWLNiW8x9niZDMDuoBhmHud4ZzlKzLHAwmI0vCNtj3nxI
Yl/nJVC+QzU/7OTbYyFTt9dlrM+K4z15xXN7pCBV9EU2/4tlWKfgFfoMc/Nn6V8NEsKEzXPGn8dq
nXczKAoeKTdEeaVd2+Twn/0C1UArCB+ieELU+rDtA/lcIKIa1gX/gft7l1b20laMPjMeMmAoojpW
RXaxrZz0efdoJe9iEeq2+L9XWhsStdiNP1L8esdtjwdvwQbUDSVhpQqZZtyePVo3XwsS9f+KP0Ho
WrNg0mMfqgkEcT+GbOBxA5tBoMb60uArQuhTIuf2hvqXah16s6I+Zbfkn91QDFjpKNzgbTTHdA/X
FbQmNMPSe/HR02+vHGUWhdY2sdBbb4l+QaAn37cQQgee6WEappBR3dbfu4dVkXLbaHeYd5wCB282
w9OmDUcBfI5E0ZyrX3raD1WRW4VyC2PcoXPtaHowvRj6ObAU6p9acnBiO90yJWG+QzrHaxQ1GPdb
S4lJPFsdlrKwTwGOcRTan6tbnhg+Z7hEuKBUa40RSXT+fJbTiLtvQtEYKziXAzZwjqUZPUQgULJ7
2DHv6utDl3XXj+54Iwofzxk7S7KIoDo2W1vBWg1zlgyuGLZvVrffFdqportIkZrJ5YKWuvV7l2rk
27SNU4s9keojdgYPSv6zarAwLC2WvkhiBAflnTrqhJ0lCu2WhM8DPRNatu6gZfrNgat6Z3D8vpkb
YcjRcqcV4KWTFxqvlbX31PfVJlzfsfmXp/cDGKfgM1yYBw5gpvjBWiKwOXZfsyuSEjO+AhKmoBaC
H1u5+V9aZs+ODDPNWAPfQWdAx7a7DNmH0azl68q7tMUEOFR2GgCtOTXCGhKrPmVn1iKQuT0neFDr
/J1Lk1vfWRbyU9lqHhl8vKwaJJr/TKZfUOGVZRd4lpVtp0xpvYX0ZOYfSvSufM5ry9usDeTlBS5S
sqa1YMGt27f9QP1JVZQdZ/G1AGZcCNUyD+jO8eyqQ6PyRv2Vpqmni0IT8e5iU45348RtVGAaFoFD
u5xM5TVE9FVE72og/eIY/4BaqiHhpwDEPMkEFbQOSoMZRdLC4uYyKJJgeqjQ7kNqkyPvVUgnNCGX
ChOZmMNRLiT1Vq2r7ZxgP3HGGPrOYCmYVO+7JlsJ9PWWyfX7p4vMjhaCoTRHRpVob7zK+8z/egzl
qg+CQAL4eZEFTRwgVB78OIuuwkX+fgDNzCGj4jrW398ryYBX+Wbl4oj2Hy2q4d41uGhyxNo2LFmY
Fh64qkaQSWOwqE7kgJMR6g1Q7aVjI/EDJkjf7vmBlUOPqv9NJWveV8CrBaoFv2/Ywja77X49PRDw
oNGH5bhO3BSqRZY1UkWgbc/8uPtBY13Hdn0l687FksE0nwDlm8CtRfgxzS+CvgcNLcPyYN1agMTb
PGluvpJYOHX9mGQHdiAFkflY7xC4VSUfncq9nPb4DngjhmACGVDhaPoxBUU3yj+COCe8AveSy45y
Be7WkfLIqB0sNR0MnQwr01B0gnUtV8ToZ+UrDliTyj4v0rn9McM/VfLPuXFgzb/HYs8uoQ11YO4/
5YqksIBGr05hCLe8kVBtSD4mUsx6TjkyoL+1esD8H/kGXLCGQgKtZC2wQg6Uf5sg2X/EDkKVkpsH
hQShCJn/kOKHcejOzAUt7RJJYBfISTl8TNc/yoaCdQiXs28xoHptHliMtIWY/yhN9g8By5sbvW6Z
aJ4n8nV4w7lMys1BCUrReK6nMYBXYIhy8auV0TO/4WHnQ7QqXpCnID94FIXrieAw5EU+IKF0e5hp
OYY+9QyiCmGtfQwg/HFl7FCfpIkSCeBAMn+xr3mE5XtRFfU1KFo3oqPI8Zib1vKljQMIX38aU82Q
YtNFjghbEZY3CcJuvZ7yen28K6YnUl5rOazW9Jtrbh8lHX11EWF6FX5QlLJV7kgEVqDEBieGis9i
O3vg0yyJ9vt2LIiWXYpBY9UUheS0jYdKcxrnG4QN+70AwFaQ2/uvV4vSTxTjkWRgM6Y2KQjXDVwN
sa2H3jLmdZP84tnRQhkT0aRUaDgBFvoE2jZioVl4oA7DadipvJh+EPQZ/3SdZ2sdUG1woPmsu5Mx
psgsPSi4U0+KJ0/jF7SB8Tq5Hx+AQMXeqnOtwUJBCdRl+WoLaGAuTITzyCxrNKwdCMMy/2sZmNvs
tgkjJOzsgH5K791YIchEg6svMaYdgTYw8B+TC/KTWiePvrgh6qKShr48AmyJgD4ErXQhZUSxVBSx
feSAv8o+0LoLQrZpCNRU3KkHSWm0y279IG2dAw2CUzilqvh+EulFRZ8ffaRFUIieZxUNAnGbgTGT
Nywsrq80I4X4iqaBl737MgYZo7tFJjA3czK4lmX7CnKXoEgWtoRt7KTUQ5eeN1w3Z/JDKGWiVGO/
kRrGGHCQ3qwaNB4MBbizgxoIJbx7OxGKsugoJIxpPO/filNC5kcT7O5B83cKBw7pO2gU3D+iIryH
gy5R9/Bwc0OgKucssc407iZnQszNx2TYAuk70jwh9kTcUAXy2h/yQefVkf0v4bhIRe6UycBR/GFE
LWmwcG7CIlU4U+jWhR3QdL5cSSNJo3pf57CyUMAosYaDb+zy3Z3EGBbXGC75lyTZqFmsgLRUqZMh
rqPYTYA3R3/cqIJFUGvzyLtWX+rUJffv0FzFMTPvv66LyvlxzBtqZus+H6cSjSBDyCnPKW+7ZdE2
Hfqp8PQJkUy4m1z9fqrF8X7tF1Z2xXFV2l0uEPt3kQB+CVh0lWwBIBJ/EO0ii9UbsDi/kyDopw8e
yhIRI8waeeu2wV2WpoEEq4N4faScPrC53soDt0L0c7jFYoHVFoMZrqVkuPJSaoI1Iw9Usw5SkIND
i56x/SfnBYKg6cJH4lvxdKxS0bdSHhH5UJYczyRt+DkEoTPPge6CEp5VcqiAAmbFYwX0atXKVLvG
Upd+WH7uT3x5LfYDwc9ZPb6iTz0CqXyjmpqZAoK2lqpN1QX4QcU+rF5ca8SMLBsbCDjkOdHMsFpY
+IYDiPRQH5yaZ377+DCv9UsNWHWmKTrS9R/Ut8mybHvfFKig/4qNMOrNmUoB3zhD6bBYt4j8TzXa
sJpv4pJJJ54A/Fokm+JuU7Mx/lF/NrmgWcEEKxKvk2c6hD1cUe/BOap4Ey7nXizYwDttPnFba7wC
f2+awVt9Ffv/u9J4iSNriEBJpP3QgMlKkYLiIpqWhTDWXDa/PNHhe4uEMAnRpLO9bS2uYE9YJx+5
0sV2tpS5BOBLLVdcY7kzW4WWlyp2DMhsLnh3KCSItCHlue1gRx0jyIGDQWSmxUYMVj90cQJR5e2F
W30l+dBnt19Sj3dz2BoC2BBZuWFs8QZTP5jcHKZ15m41DkC3VHru7IKYZ7pcPLBmpXEUdnpuTbZR
Mwcq/J5YJNuDDxsdP40JZVR+Ax69+lgxeFq2DE/pP9yBy46vtUpa2WCzsu5IRnhyqwJUV+yStKJm
NwApsQZFUEml8GmTNDjqqvOzk7Rjnz46CwZYRX4XIjKIM5IN9MS4L4Nkr/UUxh9mF8QfYfZOYFZ7
w+XeUATMfuS+RW5dc3N9e3czhxb36M3gFUxjmgBYCJT4VP6p+uk/dSvYLxPBhdKVr+SHcQtgytGT
bpHFYTj0AGKmF2axLJTpWNR4W9wc3MR0dy96S7/F30IWMdcWD27yDBYXHNdZPOoNRHaXJyW3c0L4
XxSuVBWT51XmNrboHSlYhCO2tLfebN462rutgGaps+MaWwwXkDtdv54R2eKt7wdUNQgjk+ZoR7wg
pD6UKp4hXOZNBKeauGn3urzAh9rIC9M/zBlg4zQmchVyrk5myjqNGhBXpDMr6g6HGdqGCM2QWX4O
oO3mJork7HGq/ddquu32QnJWwz74iB9BeFxmCytt5f61Ysb9i3nUOk2DD9efYdYJzaiLgz/f10Lw
oqF9EzWN1UGMJFMJGo2oUA7AuSxPUE16XmqJPsNGvXo+TQnD4f5jI9mcILBgqXut8pusaFGaTLg8
xdXkvObHh3zzuzlmkhHtV5CaN1zzC6zU8FexnVjUYXQsaQBsW+CmntC54rhGkzIYQQ7Sdcwjb7+Q
Ijw1CrFUV6iZyWcV5hqzAoM7/5/dS4WSQYhPdrlbIGv1+8XnSgiCHaYnk6hewO+0R0XkkWkV42bt
NKcKjOkzdEdVO3qZUnVk8ZSaHoDUX4dIuoa1cPd0Yc/ZTkuZ+wrbN3mBqhUoW/4wWMayLgvnkFJ5
I/yY08GNF5NSwy0mKzIrg8trXxwkcHX1jqPDfZb2MBU4AObPXvpB5UrH0x21CCBq2T1g4tNCZUtr
K+PTeHfy8uR/zdVQ8wM4PFadOO0YbgMceBDgin0GTHxarxsSYX0UM/ZvIpYNJU99CbGT+vofP6pX
xdzNyVJmAOEBZHC/Svw0kCGYKdCJHDS9zwfG4Z7x6gjWZRVesLS5VXUZbw48KDGPQp0UmtULtqzx
+RWj6VCPxYfIJhITVxm93l23ArE+m3nlDS79X7Q3vXbXgzogdrlWsCFSrzgkShPBz9l7wa0r7oCf
2rUTphyZERzmoCEC+CnLozVIeDi0RUj0G2xxYj5qDhvjxXQEqHXrR9XofqnL3O5k6Tb7Yud6PBCt
Xj5uD0wLnytd3fRdLsPCDyEqD0wQh6GvZg68eY4lagjBvNzvsZu3aAjCbgnI4XGtHzGQoaPE+Y+k
336yofK3fhJZwvr5/eQKcOWV5H4sQN0osEV66fbJFowgpYrGYl51BYXhBuWQLScJ1Sby/xiQvZbp
vbkfd8dGTN+KEBXWfUOEn2cyAnlxmTX0j8VExSy+NTrmIfZd8iSZS0DbptGYGpO/CUZkW5zEJd/l
ds1cZD5UhthPcc98QMCAqzNvAauhn9XAxRhwftmekS3E0jsZv7uujroMISLSdrts9+Wpt43xyEg9
7z2SICedACsbJBXwi2P7LMU9qf8CF7CnS0cy7dRI92MK/0FPnTvldsDZlNSYPLLWwv4xvxkxRDMA
0OthRjG/jXxn2cwgXw9+1gKq78bknDjmC7nh9lbpBRsPfPSvUbp2k+LenXYoXrpVU9a4KeAckgBi
JNV8nyeubn5BqDpzLhpG8yW1XZHfCL+uD4HO4Rfomyk7SoZNu9RsX84dw8D3d0DE5yfS1x/WDJ/z
sxPbedwffUwGU8b5C29zpZdrls+4/yDrLgO1b+WoJYM6YiiSOQr4oQ1c67FIPReqdDa1+IC7kDHb
WzQNhpWq4nxPE/K7JNFpYbIIlQgY//SjRZaFxW7ABZCGXM8vjpKgZfhEfkdi8Ryp6cEe89TDJS32
eSJY7gZ9jHUIzF9BUdUSOlxOVOAPQ/HfWuwzx1NOeAZ/u4pxirfD9U3WXyRvyHLP+Vsa4hGhJLnj
zptP2ky+/ct2XmurgeHJzL5QmDPcsMeT+lnPVv14YexVK9v0dQskZ18K5XDhc7JkmNIDqCP5pZIW
oo+ca/q9CPG/eQsKGMMR/fiyixqZYVfqVMYtZj40NHZtAE5XFKraLVITHSDB6+puEJlmmiK5ckEv
79DclDpcD5YFqqa7K4oQz/tKwgBLqfqHY0pVYhzVxD2Ek40QjBjp/+ytIp7iQyxPcRnkl+kKMNgD
SS86LgH02x2zRyoRN87I7vx2dYiXZ1cjYy0wngiFyGGqkfPIYhnyDApbAdP4nXORyRtC6WTrEHqS
d0obJbQy9eUUZ0oFk4c16YR73LKvG8NEl6buysZWz8Uh2UJ/3gD/s6avqv47JsD4BkXWwkUfx1+I
rOukXFczOvC9o6RBT9qhxrAl4X7ss09sVEwjFxqTAMI5ygGSLQlpabvgD0k959Wl7UKBNNKHJAdI
gSMCPNfXI6iAASM2sVjwmjx0dg1fkL4L6iazmwIik5tJY7kqtDhM0W1P5xNzAiLDlUXLqLYHs4cW
/xzpjXjckX/pLJNz0ZjoYdklPkokZcbi4Merl2dj9VPRUvZc8bDNOTztgUAyIIGiF8OCrUTEbanM
gLSExn2g/qc23wex4MHBT7/cx7dPmNJi/kNd0Jgg4p6r3dauKZ+ukUGzdc0VUKhjTYd73wA5OtPg
h+4IbJeMliKIzBw664NuEg334TfEy/gyZBtIAuhOg4860MVHuuRNP4dPJNUagCWVP/YxV5YLLcfq
cId2uEtCi8s5dMNQKP4lItxn0qP5k2HNmA8B2kbjyxAIVSsZyqkrH9MoRScpxQcdoMKLirl3L8eT
QXqePTedhSlDyOO1vRy5m0bfRkEGpS4yXxvvHbvEyfxmq+KBz1BdcvdJoijvTrufPhEZ5uwpdZDB
ol5GBgXMKPpALewyHEL9aFLZpg3LganqLmWBURGw9gU2gD7nj7PfFmwAeoTMY5ohMgnGknaKeAjb
db8/X32Rkluw+Lhs5IKWxdZEoQXBloR3XdxS5+O2i8LBmbpU/pQeuI0PVDgtFv4BIKR1TyBLMviA
Zf/E7se9OrLp/7PwcpYbs3M1sFkstGGEniTmbGKJeR7O5o5iuVVsJ6uXDQrbnKuzjQIpRIxv5n9Y
zvZqfujbzwe8G//Bv953x6x8NFL/FiTa+Gsdkc3/yand7fm1U0w/SfwJtFDymcsDtBvQBUmyvFPh
Jc+D9UW1pxJeS1JMxuAxWcBYrC1sDzDVqPjZiWKsi41G+UHs9twPmf+ost3nqHQQdsQrfvGMXS/g
EZSwhnJx7DcUcsU6nIUAzGclRAKS4l+m9YFVMrX3xvHh6jiEXc52S6t/td3RAgBErzXKcmyRkjpZ
CV+nkIjeJ5aTD+brkt0Um2LqqMsjI0zDFeXhAVladUF7eUbFDiU5ZJuTwlUJPxThJfHNxrKpuVGE
3/WLxco6acsOle1Jxbn45g3Rsvu6mEIDBVz1CT3afbZIbtvgUdHzEZp8B9RxsXOjbn/Boc1ZMc7D
BuJqs3GLz3jwBCq1QqNj4b8AuY1RIr6Rt4O/z7UUxRFYxmY/wVoIYcxxQD5AsCOeH5gvVQRav1rO
wShI3CJx2XvUwJtSX41TaC70EyAHUxjHNt+Lklxz74ryC4P3emXjCvX3vA3sFFN9GrDNvmYke0X5
LxdgqLQkUEzsYWZyD/iMbdRTfXWu12nhZ7Ck+shCNzF+zNAADoDKhhMZuqibN653J/klkNuOnvI8
XM9j1s1d/wNMyUQT6tYAF1ZeojbqiVyVCSJ/qpA/eJrVF/lM3aIJ2HjdkUHXs/Bz2eNA7YHJgVc8
C7dwAVEl+VZj5C/EFBWlDgrXjwO1tgjBEn81NCkMvF7d/S96SHZeeEo5aPhdPr8lqSqiRhwKEQuB
HTgoKzXir1FSnWxwEtNw+LE5XIJ/5hK2wMVhNIDEg/9xfSkRRaZRiZ/ukCFxB90M2VmnZhq4cyPm
Db4pf3mVDnjpnxTJW0ggPExIbSUupFCFb6jJwGEJ0TjBUazIbueTRlCbHIcBG2dVvIVLqwQD0IjV
H8/6IYVgD5htvU6NvmoaH0E/da+OJbDTGTML7o62cCxAElD3jJBLhX1IiIsNlaJFFphiNsVXYb0+
Q6+f1ellIwdGKe913pWop6nc+okeiw2zkUwspAVQczBwBPlCEMxwQoXK4Xl4/p3UIzkuUjhsU5YP
L0qdnN73C9vOa2u/Sa+cqIr/bTkZNLed/8mDGq5J20UoWaikWxb2v4/tmV0XyJsMg3BeiONILGoH
2noUnvUbDql7Z8G+Pw7l/xUmwG/Oay5GdePdan8ZIksVvdzMWwI9KKO1ZwQrfuF+fLu7mDaZ3lWi
jglKvGrxtN02KJnjanF+ihEYRRJ/molbCPDGKsaKYFHzASuYAZlK4OFA874ZgqhfHjRLOEUPKYfi
cN2TOG9LzTkXTjlUW5J0Js8+txpTPfweJuOUBqZhBWJBLST9j8y05JgbYMpKrSPK/wWhmE/wyx3z
SlFVHI1g7SNH1e/mln8KjGqosJrOpeHSD2ERlgXvQQzQ+0vGmq3ryD/MvGG/OC9xJTa/HB1d6Qyl
gbJKIBxJhe7IHxwDN73DzeBDgJ96wh3Qx6NpnsK72Nqn9hnABOdpGQXhKb9BQlHgjsnMiLCiZ7DL
f1M4vK8viHZEFRSVF8GMIrl8tlpEo77H3tYtZUPJ517diaVpnmVGyNfFut0eSCADvmuDreoAApWk
Zvi5GW0xJyuBLMR4n0x2yzdEaJvuRozX0FtkNxvAqaMJsErk/VizYX+wrLM7LjSpafXQa+UKHbUx
8qAohIs4EUtrdkcBqYnzvCPsxQ9ZdHIGoIJA2y/wx5hmMQ5GCT8Vo7D1Q8jZbGcPLEPwq5p3acNt
GLtX0LXfB/+65T8x1tKs9XkQZh/kH6aMyTKAgbZOpmox7FeyUsYvXL4gYKMC6z7jheK5EgbMYJPx
gi9g+DRPPiFNQJ3UnQh7z6jnb5XJl2nNnyvyp02tobD9yMXCKWzrbQXpEI1ic7yvGorQfwVryydU
3tL46smYrwKoibqUihnNwg11pPV7ZHTENMWV3ee/0zM989ZiRgXGr5TaSo7/bzUVSUHy/CaYjpbc
FfuRvPtun+sh3C91Jiqzwe2CxOhaVzJ8pv1jQIudvikAceQab/hW+7dL/eVeVkYzZEIiYJ4VKm0R
YAUhZG1J2rWGHV6ke6mBkdZ0kyLOlv+VUC12Y/jvZIlXvA7UfYmL7uItoqAw3BNFSWBea8nK3eF/
dmpBU7DkKVaAL6h6Dbkc7E5d4+G5+TS938Ih4b5Xf5xZzteWG+IgpDEOL/jyQJ0DByr/7Hyrhruz
jevUAPCiEJ3LMZR8Os/roqwIce41smzIOsjPy9rti5R+Styoiuvast1S14/yM0Wr0IKiYvK22Smh
/+F67TgipBsF87j7ru+ycGuIRhdi0sqryZafyp+/xf9oWvjxjYxfHWH0UOIbKkj83u0yVAYhcNDU
h+yfeE3/sd4TrtQLHgXbOHBiRigrbHyZEFX4Qa/56e42xgmgwXpmBiVGfVJSDeITHT7YcLt94gyU
kgv7ZtaJTfERXecF4vbF6BzhcYEGcMm0b7AdBbOcquL5JdM86qTtyjFXJ5CrMWf2QOAHlEIq0Qhd
YJvpikrQ57xTvz2eE1Agqf7D49gilXTgoyu/nOXxn6+URn5690ItrYkshMPZcqJ347ZPYte+DydG
dQFMW+gKZD65RgcbSnNjQW3YD4lUWX23CRD/lUK+heebX+bskVL1ljWd0agjXpaxDFlgXQ+Vb2sK
j6jKfUzM27ZXZ7dGy6VlTfL0GjV9W54sveC83QpKPWtNWlAcqCcA4VHglpN9QqI/IZPyYhGyKeJ1
Rzp7mynd8rLiWWIqmQBvyw+/4UxGSSAqu55nmNFQzSNW0nvUkUEiZwqdOtC5Mp3xNmTZ94evpbdR
DMOz0ipiI7Zm9C9snbYqoxAjxPW3Z6oRTwtGw+pHzoZUU1OzEeN63sFMjYOvHsUnma5GTwO50uGF
WeSu0pswwBOFgyl9k5k8yakRP/yJFR7sktD3UsZTW9bKGQaBjmbjKE5ojOXjUK+le6cYj6pU+Nci
NJydzzIiD1Mmzuzzlf/qGV61SN4YbsrK+/jtTJF6tvcrVwOKI65P3Tz2MeSyGXxe+RhT55FnBXTW
OV2TPeOC5gLRaEK2D3N6cCDg+cmuO/JFz2oyV9MLyCUud0MBRdkp80+uht2d8QLTyKSKvjT/TimZ
9DCEeSKuYhOcDpJDwH1OX4LZbXO+8Uv+Fbiv0qf8098RztWxNHbZGTRGsp//QU6Oqmc9yvNQFBqW
xV2dVmBg88yBeWvmq+mkoroAb9Uxx6EZ+6pJtBFgJkr1SHgDd65Aib5DAVWf/VIIDkAyhwsc1HGx
wKU1L5o7OLA9m/yTny7lXlJG2MrWkMkz7SdbcUvtqfD/e3ABYVQ5J2xcnhwPdOY4TKOf+UdyhSGr
xJ9VaTXjN1YEDIXxyBJmMGckKOS7hlAaPrsEF7nyQSnxpkbiVx1VbEdc5K/xbcyGPidrx/gOuMk0
t+ANE10ZJHWsfsZy7Msb5B/fKNYHUFASabdN0/65oQ7OQAOI65RcdXgmHGloO3vSkn+CdQuw/GIq
+B7cPEK63ejCcmHYfUWtbuSa8vt3Gr4Gqnj2EmXLBtmyGonlpuG4oqlpIV7+khZchJWu6l2dmBpk
/ug3EZa7D8xYPnsRqe2m1UZVuWFEqq34ZeIwaHL1dUD3odwxahVW2OsKnjyfFc2pHcSS+jQK78nd
o24vN7ydRof4k6I7qWbCtzLd5BAfigZ6MRs0DJNUEKJem1+0g/bJmRru/qrEQXpSSq+nMpfAwRgQ
Iemte7GCnuoHRYddeIVlBDTRBgmc/EzifhxxDyRybpm1r1d+Id4VzdAIseJjD9udTVB3+ghH36R6
4kG+b2+t3+mHPb3mok93r+xO4akqcCJYAtKABU1o8PP+rlOpdz+CLCKKFjAmq+kqeqm2r1rAI7SD
e8LoAa1kL/9cQDKtowgabuG4DKjXXRRCpAJyepxP9GjXBvsjCpAZgSjw3IzS2I/q1InXeuY30Oex
zUJcolHaQSGwGFb444HK3XgSL/zmSdScdbezMbETUwAbZpJA3gp95bRmJnnb9LauBc3KLbkeMEss
vMZpMUniT1pUfkqunJiYwgSQY/o5XF6PhhTxvjd2HASYFcYt6LqEDUPc3CiCBZrAd9eWabKpUr6K
nK/TR0zOnZPbu+a83lQm8xg/SjI8EF8O9s4ZfXXYPdj8BRIPv7hKKoVFU9Z2G3IUdntfYfS/9YK/
0WidQRdspgbJ31HUtj1h9mjDlxx9H4pZqGIiAGXehcVc0da+FYlFQXJs5AkdE4JFqgePhzJNBMIx
WPacQ3TLR2JGdOfsJUXc3FDnDFG1lYwSW2hv69X27ChXQDDOPFkNw/d/wgmkyaSmPi3ANuDI12Nt
EoQEy8AG5R0oSNISgThrD6FqWoNJNs512nGAdNT9znrInO3CMNQ6+OVZeGqymKX8ogKdTNyQQ6tV
mfugqjVS//+HJJkGynFSYOz0HQrgN0T8JZq3mK/Le5pjJfm4wjH88akX078AXbvRluqVNC1pGlEh
iXzZiiKJOeQ3xqy2xAx0bDSNkqiCA8mxmxHmF8ke1OW6ocSejrNupSo8YHx/QLeX1uPAUgCDpdEu
JCf2mc0EPb+EnZkiVSm8YALjQVe9yJxadPMF5ZiaSMqWHqBnAjZ69KqfHOBiI7fKSWZoIGaEwuC+
+cS7zqLlZWrH3NR9toF1AW4pXLEnJVEbjwo+iUNbstovAjiiz8DQe70QGTv8vN7/BsYXlaLc7uXE
iFmHEMBbXgrdY1xP/0QO4knah5EqcIzMWInyEdUjNhtMMn+kDEBvDZXshHpfcoBj6o5gEhemCb6T
XmGmZlr8DG29Yt2wqvougE6RuLULHYbpXZp/1gYG4cf2MYkpRk9rOEEvwUvdEJcg9MXokqLQieOp
yYQ2vHXR6WHkKHaRSK3EEdB/vf9mDUBA/kUn9LaLL5IjqiCKVgY9AOa0gYF4h3NfbITSXJxdI50H
S6E0/GFBWUcIUwLIhzbKEuz6xCNJ/f9ZCyNm5fQmNGNgGtPOMQCk6Zi9uOQ8dwMA2VNQxP/5A0U7
FDf95GGyXANQsfoYi0gEPF0zRqkwRMyDneh34qhV9/mv2l9aOEYLiptkslz1q27+wnwK8U4VdplC
s+x/OVSMSSL6Rglrul5W5jBFEzzpzQ6Bww4F8VYF/ZEyyx0qZoG6nfL2JcE4j5PGAkjKbrtVZ/5Z
mnNYBkaTrCbciRfU3vBksZIUB7tg/Pm4nqwmyKi380qYSpx2Pdkq5D1lJkWhtlfFkxgPybM1tf/n
bxv2QD3p85LC+LaM2fPilmmNnkxa9UWOWU9qURy9WozQCnoCYGNe8H40GiPNiFlNUduwqFIXfxaq
dybatLXj1nppHx+9v0l7QCzPzbsp+h9iXbPjrBfjdm44gCHZr5lTxWjTD4Fi5krP25cJI6fm2iJp
/3eR7Z1tH4darkIqWPBfyr1COCSP/ipPaw9r5qfAFFaPhJ2HIZXnnWh05AtmDVXmypmrE4IJLtgE
XRvoSDV1z5SEy9P7aM/wl9jMLTA+zPnoD3+VB2c2J/iuq6sp/g5CzF2flFf0FIwsTnCLjdIS0mHM
3X0irRstf5un3sloWcNy9l87s5UgeS9kWzcb7Fh0GZJ0a4zs86IRwC7LgWtK0kflzZ7zRXHhJP/5
df75yyAd166xJk0MmBhZgOYxJcj2qyCAd4tUBCk8uGZamcNDnQap5irmAm3mEHivBsQZgKMvGc0y
kTI6n6UGT5RwBp3QVjZ7/rZoHGOTOBFYrR0QQZ/hQNrMYWtkTt33mYcsbzdWT8JpuAQ769a34jMx
Ykk5FbjbzgRqUTW6kBqlkxbEklAXEsLEVW5/XeIvej1Hl2miO5OsjUbR/0y41OzzSu+9AamwiXoM
7kfB3NthdTicOa3QGs0e6EM2SBXVSP53+Z+/XrDCdQsCB24nKdRBKNcfCnz9tU7VsdH97y49C1YF
s+d+4GgS0Gu2cHe2c8EvuOBgdKBAXV87vBG8oVcSojpmASBQ0GLPiElG8Kxj9pgC03dwW6k3kWip
asnO/chMNhQvSzRKVblPx/v+YzWAK8gJvji4kyB3OpIiM53f1CtavzSSpSBusrryDZ4lJW/g6v6o
ZIfZCNQecywpv+lJv+mFdi6TA8WlnrihIXfuIr7o2yYAj+QPnz/K3ISB0XHzbXuSJO5W4e6fFsxz
VRiaw/TdKjtIdpNt/Z5wXflYimwibuQAwxz+15MPGuF46FqqCycdUYFqMJK8RC/C+OroR+Nr5cmB
825YtNr/yc0i+Z82hoEa6GX42Jzn9LrzF9gyuCz5a2ab4PdDXtpyYJOSocIzBFMl93sD/LItZ857
CLxrGEXKqP+8kMimzOgzP6oi4BW+q0LzCshI9x6HmGyjAmpeQIyqMGmCxPi+419bpeoSr5JI3RgF
MfGE4GmsjwMMcCjo7hxzSIzOErSzq7QFtdhHY/M95wyeDGgxhWLitVMa+A8GgP3iUuF6RpBHM7pv
uOC0djWpPtz3u/eYsi9lZLvrpFVoUyvzwKoVcC+MERGrkUlcr5EHPql65yDzBY5Tjv4lEYTXCgVG
jM/aIJ1GGqaDlL1IukNhR1Gi9+pQq52GaE8RFR/SykKhWYtTwTwpEE2/bO/AtHieUiQ/tvH7pySn
8Fmlmrk/ihbMT2QyAYThsVe34Ebl1AnIYWLYQpLaz9Sm8gStijnwZwyh/G0PtvT2y7/rp9dfhQtU
3D/pQS5cuFvBNw+9WKf3z1boJkdO/9qePPvfUg9lrbLBFibUrbbvESRm6uQ8PZQD3uiHbZ84OJwA
zzrejnu8DckBKOMV8OkpLlfUjLzC3NAwJuWtTkJjqXM6++OXAhJBYJIYEcka5+nt5JymJ2BGlj9S
MjjFOjipp73Y+TYaPap1CT9Cf3qejU0GVuPA/WpuASI2q14nCe9EAZj8d3iLnS7OXaz3SurmlOAh
QBcgpXYCkgMc8QfoEIEba7358cR9Ot6noVAieDyJGsojVIpOfxXFhMwaSmqLtngwJCbopX36A5Gc
nUcGAitdYWo4bFmjhgxHKwWHc8Z2Eik24VO2kgqDsllzEt55Iy0x2QwenJbSzwKMh91fL77rv6TU
z+ALPOBy/f69x4Mkd9etYzCNInSSFY2I7CFP1pIkbJx4u/hdtkJO16abn33ID2GTljTzvR9R/sN+
0DCIQFrL50uJuFelPayrFh/atGiW8YkBwt2z3nUTNxKnVScldiujFvUu9H9QJcctxT/VV59M1bHp
cBczlGKwNwA8WiLnbuS0rcQjK2Jmf8ebd1sczT6O/dCst8dVKDBOvaYP8ww5r+p1YXxbyz9XCd8J
b24HQJ9cfZ7D7gLNMcjVjFltkQKY+9poYQ4dhVEKeEj+9Ur0PhrmjOQOJm3gJgqhgLPpR787vB23
bVioFbVip2t9tkhNCShMmeMT1GZ7sFSSN7eMis96RHe9GB7Jb5BfsCC4lVvFYEJ/KuDtv3UmtBCq
h5Yb4gMjSITok65nKV99i4oxynj874fhSvxyuik/BP8L/JX/fP4DKd5tuPiRhPbk9BjGfWONxkLx
8RReZP/hmOalvuN93oWKljiyoSYpGk6Fl0lnI8aQF8HrQaTlJSEW3X+bCLxQ9DLeAkxTctMdAiAQ
OWkT3++wAma5MPLP084oTep8fMV4wKKdwuZ4QiK/0VYw4LciZ4XolBvSUNl29LOq6WbeygjIhbe/
k+eEZcfzP37nxoiyLt5Al5Q83uK40tJBDvFEOI66/lQmhskRJCBZre9JpT6b9IH8evG01wQjlDNY
BNHikxvifsRotSgv/by/Uz6KUQJFDFX9OP7QwUiilNoSR1qG+pIYCtJZYk+MD6/NTHBfnpVxAVva
jKRm8dTAcogBZq8NnlMaRETjpwojNdOKCPBEy4y1WlV5nsz06K524pw7RUNoCQaSKtx0CPoicLgQ
OlinHADt0tA1qwKnVswzonDoJMDdOPWkaUB6uqKMMbpfT3GvSQTpe9v/k5dq05yAtbxuhAWjRZtF
ZHPbZB4SMEfo3RZ2CJtTbWfl2VKg55u+aD4rFXr8kE8fI4nxQv5S0KA+Zni291L49XsrtXUOCGYy
xtOUltGdG0ZsO87G6SMDCqzVn4h8ReQVItyN088Tnlc0eMcjenLn0HzkRkMZkEi/j6YPy7MhQGTh
+pxeocwGEwNk7sVay7xE8WPJhM7KZ/tpCdJwT5c9uxMffiYdjUwr9RYDhycPqxsMFKYkgw5q6giA
wKHNNbJLqLmuW6p0nTDvsvMILISRqQkaUSRVwMRdf4hRivQ+IWwJfoseKqlZBvqV9iXw3GthsGUz
xJ8jDe7efrzJNLoZyQiXzEGn/5CIOUiDnhJT9u7JV0adcF8Bf4xe487icrIeUZde+IJz+kijx4k2
ivwo3WwX+nRrW1ejC6s4Q862Bt6WjQJ+mD5Ax+9bIGF8/1nazAEcghybcuvUF9B9BlziZEKT2l83
SzUzWakSdbhghPK5o8G166rptgZOlGQwtKNVmVubCoZbmLwWEmkT+8Hc+l7FC1t2AWzw0yRAvcV+
T7sVSodaRIFMC4RX7B56FpcXMFXKlofnMZoVbw13E3bIwAFtMTVTuw2D1j4lF92wk3GJ1OrjXziI
n500VXW7sFd4VLnfzo3o2EfHEbq7iSkeW6u5xpAaf1yuopc4WqOs41JpHO94/nEJXNg8tej+NclT
hYbRDA09ozOg8N0CS6ly2bgkLsgCrKuN8xQQlfrxNHwafnYN8wyRSnOjSPQ4uecseXUqVCZMQjeP
laMae2xyEqm1xtrB6K/+Mg2aIOm4+OIcNhZgVEcAPW8U5C47dCbzzlNUk4DpfDd3YCcy9omwv6NL
8ts9+o0ZPAB6DJNJnazq1Z4yR60M2FQky1qLRQ//exRwdYe2T6dGCwacjGgyoWQD4ZRjA9ZtczwG
0S3GqN4y5G0V14dt9wOqokST2VKN25dpYaH4u9sc+bkXBgoCZXthU3LzmhcQfcKqqJtOtaTyKva4
8w53v/ZUJ2Skmk0CCB2+g4BmOoRLfXPqK33ulOlpVPZ11qGl8ujxYhhKHwQqyH2npSOantleGoxk
yLoDo7cOUoSXd/qX2MxY4+tzRAsuig9ZFJWIyuFp/bD2NNaaRyLF2ndcxU3Z/umNjHzwtcQhh9ko
4780QoZvoiGZCWtnnx1nxDMcysoQReJ9/gjPtHNr3j+PpSi9PiR/VvjG8LJRoaP6+5wYu4YTOWR4
lzUh8KQQ6doapkW73Lb8WK6309YXHbLExZkv+ZQr8G7/+G1AYzglycU+axLJD5a1lnHXQk07v1aw
psPstcHlF3Om0fzEGqI5dzj38Sur4gw/4m9kDUhZawPSKX600WEqflLNYty4V4/+utJz0UqGsP2r
jbzD/O4TCa+HsSIhEgVZt8X5moah0oIsxZ7OffS+GAqG9EAkJvKjB7plk/6rhfj5bxDPeLt6BAvT
1Wvew1zb7lRBWnt2tIY90SxFOUifj/PEaRKcTFbSQT0Wk9dh18wStuiG1lNfHxiS2ByfRfC7imRu
uhBnXvbYRWs5syCV5Kii2+mzI6nypJM40udTknze57AgW9T3m6EM9a+Ah36FxY2bBn7GrxazSzlx
osmz+qnNd+iYgipDs+iydqWpdPsNcdo7uwKHieEkdnLql9L5Em4n0A4XwtlGXISif0l6XoQFw4B8
9tejCRVQ8zbtx+ui4WtcPWrfot+87m0oCFSc7hfVN6LQiZ/EG6vs3qHR/9bwtXjbreVZg+yEaBb8
ZSX2gy/JZJ7cldvHixXmKDuY+D1WhrWdGT59hi44lciC0Au7WlJ12kYVttRouYxDMiEcJvpkOKUK
yRv3noCaKWmNbfTmyvGMlZtx7IHxcwMKY8WVMPhWcyOQGfvMIs2+KL1Kz/gnKmzPlWnXrQ93PuKz
Sx65ewQp38bC/uPZc0/dswBazRNXe1Rdc0KNA96j6I+RJHeSwvljO5CfuQnQjUl5fEt435CMkrrt
kT9qIogEC41siIRmzfX6qC4rKIARkR3Fu/S90LJLpp7gL0DG7tKSDI9VQUNKSlvw+nkSifHG9m+t
XNw69okMFefXTY7UgRyXJjm3A8CptKampkCpe5M+lSm8YI79g1c2ncOBIdQCl0xXJt98ez6hx23o
I6O+CHQj3EYnssN6DPmsWzaYQCC08z3bw/46FF0ftDOaenF2SEC6t96ks240UL+JIJFmcztxmRRL
HH4Woayja1+9+dWB6HQ+D5xa7AmHVn7k++Ip27S0EJmfIs067et4s09tL04moss+jLlMRuSbxzep
3CJu2h/m3PNlOVvga+6x7KwdwVBgJsdDPwVNGM8diNwGE9NraFUyVaZpuh9NUBVgTpxOubZxc8Au
djMAg46cqa34eqSqSOHg+V/5hBu7tXi4odO2J0Ec+KxKRh3m/R1o50P8LybcV1iM9pMlh7/P5vGK
GUn+Y/zSpb2HJ8Zw2Cz9ytKgL+edJwzAtq2PqUaAOEYbtGolPqENjdnMtYH7twbSBGhlsDX/2cYP
H83V4E/I6p9Ca1EKlQ8A++J4wpYrZPdC89SHOjb0dEgGsqwIUN7DQ5aTY8w+w9WZi/DWfiWsIdAH
9CMb0KpKQd0xeiJdUH+jTYfCKtYhG8SHpkyu6GKKgGMpIq6x1aM+is4b/HV386QuXTZ8ZsJX5JRb
K6ZOQPBEnIhwqMJWTmGZ5/8mIiFE+bYBmdt6vqV0703/3KrQXf3el47aNWS+O5BTD7mwXZdfbVvX
ZTIw8tSjujo4jiXKGDdQREZVswzdvTawVZoJ7V0bn5vNy+ECJFmEI0gLITN+Wgr0SOuZXaVTLuz2
NmFqmSfZsps6biZwyybuLgzlSTmfnCeL6TypUdUFllbwv+Trg8MNb2l2Vw0iM/BsTa4W1Lc+0+hU
uSsRj4hySSop2mID3gmDlhH771c5lWrnG5MffaAwW6N+y4OQSouQr5bZXcOW/rfl4nNabSfIXxwJ
NLW3mc7caJUCNBN2aE8+0t5OM//WjpmSOzeWlkLsMENHU5vSqZO5X388KoKzTJ7OFAFELTDxjAWk
DxW+sSX7ePkLja0V2n5NYERyg4YFFhxlMYQQMW6xiNgRNNMEBukdCnuNbtH/7T59SDItFCJKl5Uh
+0AC2WYo13q7ihwfZjkGlGvYVZZ20d0seT/XKFZZ661USAzB6ZZDpwTA/hx58fQ8C7GX9tctVINF
BDf9hu2S3V153rhvGlNLX+shMlKhA+TWtafQ9ojAZF2o2Dg0BDLRGoANCJmtLA2w6cX8NhYVPmpI
oKEmcng4DlaDSNZ5KKRknAj0RaFzr0/sB3wgHwpTeZ0vMemIyxFQZErM4GU5mkHUhfTn4E470G3M
7Iq3a9xaIQQf+I63BpJXJ3hcvsn4G+3iAkZklpj2uZCtCxMqVpQEFgDv2am077Pik28G8CCkK6Vy
Nbe5OYRED+n/dsGeWIX3Z6ApP+v8IrJEVk8plpWVdo6YR6xPiwKrAeySjDXvISCnpox2aSN3nDUm
TSAcZOsuwsx0B4BvdCbWwohWJHDcnS/h+n+W72Zqoe4u0KjwWozNRf1kNXBRiCpk+KSxGwmrDIox
CJkuKpikaIZGX1nuoVF82Hkdod8Iw5/L9kMCJt5uTyo7geMmGw343wl9DR43xTN4YB8BzJXV/0MG
rHNS2oRyXUYnXrdb9TnL7J5XjgQxDdEmvctvsil2g+m64f/TmKs9O9101/iyW8ugK2mXKum4130T
s6TfPjlmIMgGoF/KtaIfcRYZpwxXYX5uVAbat6roBvhb+CRagfVUhCuOtCrkqOKbgl7vAg2h1/2U
qxaIL8TcFV61/ZNIG4Nse0yXf/UrCdDrBr7vW4jaNkr3AJQs56mwBnGz6R3JEjDFYQfVuPnnmHx9
kw2GA9a9+odp0PYVcBtbWPJ/JNpRHXYjgsF4AoC6ysyBhrgmRI7/zGgu6ZQPVBi9ZsxopR5ylAsv
PxyU0pycp7iG+14U0c+neVRojoS4LrUJtgSIvCfk9O9qq0EAk6waiLJlRs6J3e+5THPoM/CeZY2+
toZhrO03CKpOg/st2glYaY5s/yuGTaK3scrXRiP0QIXfksBNLNPQnMvjUd4SzrxB24kG8rnQ8Oy2
3jtM3Xe0bAHPBgBLUSxuJ/gaHB1Fyex7OdjqhdC3m11/zdMvJjtbiKzxmh2D/WdKCMRuYBCB+yDR
/AQwcdToOKpUt/vvFj3+gIsqBVk7YZE4Jd/LFLr/PAC4bHticyNnxO+mo3qs28GwQQNgYFrhZNNq
6+TK5xU+UAk/n0X2fGr1wvgrrNZqf+C0FI4i7+M08mxm6aSdp55YjSooOw5zOcdvbmXUAiVYmHvz
4n+jVDJvceQik4s2dkToNaGkhbHrbIjuvySl+Wb1/NXZ5CqMf94eDmIrjxRZjbJJ+wXizOWDtbqV
BdgA0WVxc6oVa28VNToKUy8ymHiGt5nbg9eQQ2ldKNnU+Itxmz7WYzkeJd3yvAqINby3tFWkF2ns
ymDdylDQ2E9Q86H1O18OtXTpcQHU+0hVibujLwHzlhL9yrTwVBtowhzwZYpAhXviMfl4RW2H5W7c
bv51Ss/of/bRd4EGfKUFgovtYdi3IVgsGpnxmewUjYN/DqSBh0HLRdn86UYEssqkjXsCwaR07a1V
yEmrN7IzS7T6qxBobMxIwraM0K81GA39hJYTmnj2Jc0lswJg/TqetBKS96ztLhNauGSKP/zFlVlk
lv2mGZAc3dvpz8GJszipzgHg2rV2VOT82XX97SGyIghhNwZ1zW3/JZId0FEluqoxJbrPNn7d3xdt
HYD6NGG34Xjl5uv5iJkQH7ZqZtfiv7bS2jiiTQcL6wj3OVwJn0mPqdc2vIxd1m4DadRBYaAAtl5U
P0YbxuDivDQQEeJbFULMTbX3/SaXyh3W3XCREURI7pMazBmtDpBnuysY1QIkUMsGoWd4pUOUidGt
YsNIlYpvPNxFGsX8CCz7kYTPjxryvxdkRdhl8qgGF2Q0oyg5Heis84eSjMw9YlJrMzZ9airqb+xL
3bmCCun6/2EPnOJFtwyMBHIzXImBM3tw87H6oCnXFpJztD009mdlXVT9EgTkiCNA1qLh8lJtYMGz
+MBwycAXeWCXAHZ8ZBts6Ekzf2+9TJHeiQefAFa8ps3Ax59NDhTC8GWYHBkTIXLMz0eCf+CDOWzD
TLZjQ02TCv4xCkR1DKSDx/4tSVysZl3zAs6baSFeFTjYmJpd2KVJbL54qJT1awQWv7aU2FWtQZV0
twcfeuOyXA+4RIphDevKT/Hg0QPp37g1D/cztySvxDTLC0ViWHEo0EWgQCaVTbxqJpExwhffsNwU
V01xmX9AayMjYIr6xK1Gqw7cXuCUsNh+k36qvcHfJOszgp2W1dE0z+P6oOonqjrabMXdzQBJWjw9
wAy6DpOBM5646Tb/f378reY3MCp6Xbz04MYcbLttIZ+TarBa9350LxxmOz5BsPBdvMPmCxrPldGd
Bewa3IiPW9AXn1guWSvvK1DCQiB/Yxy/QYTch4LIhEn3MhBz+TXX1TcFAOoxjhaFUB4jctLpRNSz
vzvfTCAoHHcdvqWYir8s4G83AK0hgC0+oI6XJC1UgqcRke03bOok39eMnuEvxBVV2GIa5kLAiwHh
agqsx0CcMfxTQDj9rQZLzjv7fXGROfPVnxbeP+6ZF8G/H+xHWZHluuDg1s+LDhjYhrMGKD5dMwoF
lRONqz/R78bc0nNaOZ9kZ+rn/hVVZ+aOG3nTHok7nxLJktL0Iy1Ljptq9Mo5vojOJEOnyt2SUfq4
JRQ0S80bagg4ktCgscJUgVzfQVnTbfMGDfCcrtvDXBJeMmsiK53weBhf9FosGrAX28Q4oxfvyV+7
06WYTlWY7o/vpViciXoiYxlqwkLNQQBsCyGhNjfJrW/x/HK0VwHECs8ZxZwVov6MIYXKbuhpdYol
/8edZZxPM/cZRUQE+uEDBhG4mAY/qvcanhaM+V6dfP+oKnKgbjeekrsQgN07XZe94Qn9uOntKqDA
/Z7iIROelBxKgigQBIqz2cfsopnzrhf6NsbYf/WOPKb6q67il/0rZtd6SFndAVqopDIf5p6zTD7G
MSOd9h5LAUsTWVPn1DH4Tv04iI75YhrlviECaYF7vXj4fjtQ8jNhXqOt9SWJ0cJDMkaYmN/E8OQM
2fct7YVthYb5UgxoxBsffnBVnBmQAAmmoTCheN/yq5pw0eepdXamHDv4J+MtzEXL+43gMTsT1afN
DClQhv3J8DDYUlU8qxR3cWpTC5p+c8PzJ/NAI/AeMDULCAHRPDavEduQhxlmGenSD/anPxC2l8tK
R2Df6ZgTWbJO/300MrwtofPixzXoePKSu5oBskYuuLeeEJKX6da37T4utn8VGnJ2MOkMU8u9V61c
WZ4B+8LGmBwJzIrhsJDMf0bZ2EHXLECJlY0iQtBLiinPmzsuxZpkNBwJrr8vStVAWcv2CIFmIBSw
P1inFzsayE/WBtsUsppDH3Vr+n+vdGKtNaiWp9ZYD9Rz88bFiXCikmi7MI39U2NFDu0W1YVbwleW
Z+eddJhkGWC9EWzw+rvuAsnTHbLVxccRFr3HVn+QdZ6aIcrLqLme7HpxtapTZLp8sU+ke6asbxlK
3XE4efTfqLLNVpSU5Z4TRyFG1G82LvCJBS6gBMvsQ5CjG78ebZooaB6aUaRWRuqzrdUnuBzZj85n
wVb0XNze4r1uia9NzVtCeNCXRvPbEauBgug4W9v+qVvxPKfyFKFgvyUg3I64Gu1NmWuvNJ0U2qtU
Jyn9hC/xGUldJXwZuvhkWb5NBaIKLJEZY+QDQYFcWF3i1F4rrRgtuX+EtvARsuTCAHctZn3B1x+b
Y0J2+GzL4+w3F6InyDIsAoEK/6mEiAF/d7DHStzEpmcJvzEt8d4sroQh5WcmE4yLEz/A9Aa802B2
21ZJ4GsG7LkkRqUrFWn8+eInSsFgQEsl0K1Y8mlAIRWAyH6jTfD1rWIxduoKQZgKNPRFbvQ14Zxm
OgGO2F9T2zz86jIUJ2Hklaotwl2Rgzr+f/UMOZOCUgTk6zQ6EcSmBKRpxm/rIWnWZNG8GQMYpfaL
G1hVWFwo1juK9VNEZnBbYFe2KdkGHHRSriy78M6D46nec+zWWBJlXfpkINelfaOShWwhznrH2asG
g3PtU2dY4EoeO9+OU/fcoulLXij4LH7Kjc1VDrmHgjA2HeyJ7kuVI5Kdfic4+9nT9kzDaTRfAl9j
RdUmAlhWk3JV1o28vnLwuRZiOns72nyrNK10kwDpJGgedN4d13518JoBr9rwmp2oG/hmMich8KyK
EgVECczxS7kQGOdlaFCmROqKX2obcN9/q1DGxpb+lFqlBqYRnepTwPaGrMXSoR/pkzZBcAFnd6d5
KZMhcSizA8CN1L5YGvSUSW8qPczx1Sn+Wv/1omNMWwgQC/XuAXxlxFaE67CxB7VZMZXq8xxtc9XZ
iF5dMzpTM2VFXUfcIZfG74+YbdER1B7mjEY/tSGXfzyeUy3FxAwDJjJmC/twMirx6++yuyYrMtMO
MAArX+JVADjCZb7UzyXROGbj+VMxGh2xwBYZYgCw/7EBtTlzvllz5ZLhN3jjhjnSI7tCyc/Zz3hX
ROwQzk7rmnxp9ggB3TsJhz6remSuYw02N+HU67wSccIoIl+2/ttN70y/3oxn9bi0HIhmhaL86msN
Oel6u0jOuTP1Ox+63PRvldn/tlnaX6SNpvYDcn2VGr5vgGPNpRJ7X+vFe2sGbLN8l3oGXzU8G2ak
riLi0ESPF8l0REfnUWSbjtCgFvmGDDjYUf3F3iz9TeYIn4s9hBOZiVKiaSWGCBODvFuaYU8Ic2uO
npoASiRAHXedFBwQpJ8eK5xphCVe5ZHrD5ARplx83fVaiHxjdeMcIfylMKL8pcPaRMFuXVHGmpcD
U4bE5BL56ZqrdkLIPchE3dvKff+yBCP4lIhVXMSxIj/bef/n17LjHnd5xPti6P8XWcbwD+jADrII
DVKKF2+DckvRSpwEvCPg4OseuqDePOqjcNOpS5KGtIgWzNKgE1o2lt2aIFI8XbCIHtF9x9v95HbP
y6VFihY6H/71+Sn528IrMdu9F+YVzibfKyx0dIklmzICr0FTtm9YLHRMYCjM3s+6dCFRN0Xts+v9
S8j/KQEwl91SL6qcOOuYuYbvuV2eKo6zqAPmMG3zc1ynGfo83VZ2DPXFjjFQJR1RaQbqM77B+Nmd
nxyOHRURv41xBiWOv0oOOrg3nyZWJ/9rzfuYYwYUSJ8vdHxbvHNgXu1HXW6C51ogLLAzVuLBsUOV
QJfK9GXdQWJ+gb+IBuDzQkQo1KG7O8sn0LKsf3FDUtfxW5bl71T4xCQbKUWc37vqAfn3rKRq5uon
29E9AFJOCMQUoDPDcOMMiXNfiILtUsn2bBZsQL9EUTQRkxBiMoOefK0rTQg0nKpJbA822vX0O/Wj
qXEvMOql7ThWUlyDO77Ryf74jO2NpBOEtwNoyLmcMN5hMPf5D2IkmYCBW8cJvepS8s5uiVj56rUu
1amkp7J7BY47OIjh0x/NoynKO+rgntGr7aMfX2eXh7TWiQaNbG3+t6SFwD0POpNm9PJEP6Kv6R/5
nRgQFaUbmEhU9A/UF1uOf04XhokyZCcHNzXi8eZft5Sc328xpq2YROqjRqbYQ1LcShORhp7nb3pQ
1j1QzI80NCzSJU9wVpUFiD4+eHIa4tHczSx6IjoIPu8w3kuzcCwfY3Jtgv11pWqjBqkDN1a99B8R
ztJulk1eQn2bRfOfu0vQDuxgMG5sHC9bcyUlKsNvXd4V59BUPWhZf+E+JbU+TOjvzbkLJ5WDzDhh
qOPmlVERziJjh7rCX9QCYBkgbwf32TGLZZl9rZEGUdABsfCtx8BjTnHfJvt9NaFEYd5fGrNeit2Z
+N0k+tPHckvtVjtPCygjqcSiqtdUtfutQSkFhx19O9cTS0yIRyc/oRUCBYCb4ux/iFWHhjYHCpDk
6gCO5l0gQPMedoPQ2mw8dr/hg8sTceW++GFjb2Y4Pyn5Qa0qOSmliFMzwYqeszr0gvVGSnXlkgPZ
cCyvjixz81HCfsh3RUsoZlPxNoiWslOrSGPmIiOX/RH05G5w7a7anpmBRBriavokGg1CvdxVGCXE
NNrvq8+H6V1P0AnJcMr8E3AnLOPCPClubwMuO7SPVy+cqZ2wnecY1fu1+kipqJT1vNBC9pUiB6KK
T7BV9EBw5p6PuQPEqajBvCmfhH4nRptwl2Q7TAN5sv55cTVtzaKo5KN82NUWulVzMKB0YBSpqXYG
oN5gcIkZm/GIar6dE5idDruA7QwOlio7xXfKblEw65cQrGX1WLH+RL3iL0o78NZ9N8l2OX84G3n7
xOOPVB2pj8VaoVW6h/4yuwOaWHyx/x6/bnQjcks3nRgiuVBYIV2T+cThTC/AWbsteQVSiAEABrp2
p2mLcxdvVGTTvKPSnkbmC9We98v073Rutu7b8Q0U+vjqPP5buo/fEJXmO8xn7fYYvP4EaJSwGwIF
JxSXf7w/XbvUOQV4Q0zzOhN1GifKEMZZV/3OlSZ5bHDt9ql8Wa7kqhnA0r+eFFS2UXxhyEh/6e2L
h8kakfm17/uHPi7jnB51iZkQ52I7/xV6/itY4FQ1VR/YPOJSJtcNRVwTS+J8BUpL1Rw4CaI/fOd4
sCVY3y1OgaYpNp24/5VPncmFSY03AkP3LiVxQN9ox8knRRuuesbQ18KXsZUVfmNGX1LGmCFfNQRC
f6hyAU1fxkNA01lSo5UXTpbopcf5w2SZE0tXS3sKZrLNNmmdKXsJOOZAGlmRUwIQVC9fIkT0MRMA
5gc+UKUOpFKaoirByH7M9CF77qb0jvWW4ZzWuYigID/O96fkQF94L0KoZXR6nXkCgDhJnTci1WOd
o490po9An0oK+AUEAhKGHGVf6wkPrNsPn6i853ruz97R/at6u835GugIJxGAKUOqvCvue9U00fSN
tv1hdv0b9fbe0YGC+lltn5cWTzt4vFUTfhZohfRiVMEJ/wgmji1eLVuqKSVCSGrzp/XmXwhppjWn
ZzIzHgcdJQxi4n1r3utKKnMKLXtYkjicfaVCRxhGpB7P438uLDzZJ2JcZ1vo5eFgnAWZqyXKyrmQ
zdCaXOxSF2Ahnch9EboVH3EiiiMDkgqeE0uNASriEVZpZcTmWnIk8IYYOkVT9OLOF6nhZ3wYnvrU
D5uyurmuSG+MM4N3SDTC88uS4GMrgsMdi+Fz6Wp6vFKxNSU/agwvENHAn7x7BB63qT3jaGfi9Os0
+2EZvFyakAShNvaueLr+IwBc+fZ0/vhs0vYisQxrNmrTks6I2LyehNZxujsUwFWVf5eLXKjPFsMo
8KcmiZAmPDe1WkGcjTtl69iHFaZhCCexQzj00fqPfoIuvKcL1POeXi81Pyy9YubC0ffdY7mqnaC3
6u6ynQTz7roxzn2M9qsnc5LEvbSY4A1Q2mlSAceq2yT1GCgB30Npa1YynF9sSTBd/2q0xmXWCQuX
eXltdns0EoHQNaJHNCbZSbGvwEIiZT4h0iEZ9/iAP2elZuVG25RaCGssFAATrpG/F6uRkuocH9JT
XaCfK14p+wwcZ+3R8OO9/Ibu0NOuEmibqN8DeSHuCePwP7GLxbzHjDZzrt6G3LWe60MawaOkevym
bdbh3whyeU6n2Fkgrj86L4FxMx0dTJ3P6Edyk9yiwiv5pZH2OKR/lzcfryEZlmhSQ7EHIInfg8nj
lwppvCVcSxz0SCa/2QSNXUItSQoK5oKwrnqzAAgKpFz5qg0KGlul1MlClpbbdTmgzYD8moad5DZh
ZtsvBReXcGRj0ZZYBVUIoY3PgQJSlM+/iwR/+iF1oTGFPZoRBwhANCeZ19k7cfH6dwvd3YKcfsVr
BjZBtgqEGcKecUvhsvTUE5oHwXWQA6ORYpx51tiacX6nok7rTbRI430T7XZJBmU0hkPzwQCx+mUh
sdOCd67To1veoH/xZSendJJIPDf/GvD9MG05II/VxlwtUriQUeu+CjHW8TTrqZP10ZGlkBA2+2OG
PL1M3h3stOvKudpYGlerD5Cp9y6r9gFuDxHhAl6dVb2RJrRT2DGK+4CbvOwBQ4LHePJdj4MLaG0V
hqOmAHMZeuQIIt+B2uSolMwOfXPcGji9k+E7rpa9U3VmcJPOueh2bPhferZhF2XC+HGV9UzEmrWv
k/jrWyq1mpL711LUkxaJa6XW9gSibBs8h8WFc9hNHH9MsZ0+/l8sLxbeaUEOwQVj6HvASM1pd1XG
fnAbiIwi0RuWRUF6hhRExXF0EI1AQJzFqnwhmrvpYb0AhDs1wtNbHZ5vRUZ5qEtdl+cdyPI7Bw//
270mPFtMMJsMby804mbloYdWgUQjNcyJOo8cowPoZ3N8WgJsswkCkU/aWRLQEgmCc8BktElCchcc
4mxaiz1GTqspFnabxM2c3OFIlbjnHHEc2XGpXd0aoIHssPcLQ7kt+NSmK3IJ70RycBFkOtIKLXx4
m7aXynLydHcdrXmYOYvAQ0SAGthmJ+kp1isLoiHB8jVnx+BhZt/gBrg/toAyBVVAmvEBs3mxFmpr
dpd/BodaF40hcBfOY96JUjSM3BlwM6MNy9sp/goAkRLMOHvLY2Cs8g7yOjTTVdFvhPZyd/JVGMY3
YIwBlCKLWH6uxwnXnhRJyiNndP2d3CJkGi7D8xasQ9621F0mW2GxD00uGitl/DUVddiDmxxmGWOR
ZkrqD6z1Mxo9NaMQ2VO0p4NZ4qiezNSXEniQL9SPrwUQjvvIl/n+opYqEIWwEyXfKhb6jjJv+S46
dGhp9mBgpYD3LibVKCR3eHyKRqujCdlXFOrctUIyZE0CP+3WXsJqIAuOrFPedIfVolyO++4OvAgZ
RYtXrxyph0VroNh/MYkyl4f8UUN/x3DGE/dUrzv9gOt9AABEudilyim28xUKHLVqv+DUMGgzZgsH
q/2Hzb1jye5PjMPDMrgzieyFqWF8jCGcN8TiGOoVr4su7j9LhTlQweZ9F35BRbP8XT4M3UUFv+xp
Fus3bWFHQJfueU3rBFXG/MDtOvnPkIcbYoGI0HaLWgT1rXCE/Z2nb40mza8a4fUpsgdeU/coGXOS
GFdwxwUYO6yS0KfLy6ibP2XY29bb3KkJQl3g0UcLxMTQVTBe7GV0+waDMzYLbC6mn826JXCp03wQ
5dLrtnC6/P7Faf/9WyB4wKl6M/0ogBpjUIwMyzaZY8M0r3tQiMrm7Iczh3CVeCLnATyZjX4da64l
8IZlov0FyGifqlN/Og600gW93j8+Gvp/gHfQKlOC9wKEb9AQiGoxkPpdq/jkLavt6+fjurE99WSj
e1xIlv9efOcAdaYMu8vCFE5pgP8g+xdtqd3OYpKWXDeaCSvWk4+cHwWN/aSUD3rEDPPP37ymQqWe
yEw7HlJ6e1o1/sP97MjDbrvCRL5d0r+OGY/z7dMuIEeAh/zEHbMy40zD6rW6mR9SyosVTF0MdIan
h3eFtlrbMInBSVW8+XdE6OfxwPUfTKvcy8RGt3Q8fpdH8wQwDByQe4NOouCzjVgC1AO+S7x2SpfK
k3bpJkiBV6EUgN/0aOsIEwC5a9HJ1iAn5Gi0FidhGirWT0AbFvX15h9fp4IFxMtB35RW7S3f4SfW
UuzL1we+7pVK2zCoLF3jylYhra4X52hnTDXeISwSd4eS5mLhq9blTjLVZEGUR0TU7eEzCGzAxcU9
gAU57rC+NhGdMHdZf755ea/Kx+kXY/vp9WIhZSvdAULVxcj0ii1+IRCSghFOW1bcf7q/Jf//soQk
DP0Q4OmfBvWaNRwOYqnvQBr4pOBsN1oEiH8vjAJRqzFXJVMrs1qiPZjwidxg0jyMh5kJcQZhqCc5
xvX6RYv6UfVjKD6JRzpY/GUnFtejBMobP7FEp0verqlclfgvjfU+en0vBNdJBStKuRYmuMXytXDm
XsQm0yY2WTsNPOfOYm8wKweymOWaV4ctoVzSRm3ZyaF21VdE2HKjKBzoz7NdnQF5C5fg8j+ryZ2q
vrgOO07QMrH4W8N4AimRLeEZcSk32lZMRRTBCIzLdg1DCyXU4rb4PqfoiqgJpNW+21jKLa93AWo+
BFDGh/8DZzKzA0EcZ4Gw5jzf1Z+tfnP+2bnIaxBnx7r0pYPwD59rpsWxkwmxnLh8lY9S0aC0wJvw
V56qkidUR018WVgw0wgg0MlVc5Fjq1Ay8yiPzIhOcDE1tmknjEt/OZ0ZRwSswXYFXhFKjD1XeRSr
am0KrvDLrDymkXoMZs7zZiZ8OkuBnFf6kNux1ZQT8A+NZXwpJ2L2q3cJHbUS6DDuutwH4CJckdVY
NArSLTYaHaSkarY7kJSh+hYjCVu7y7ZLT9Eqpy97J4kFHXEAvKXkTTt2PJHbsnr4MYV/yratY/Hn
DYSja7w8NA8/Np0D8VI0vXnq7gktLFAfi2G6QHxEjTuoGlZCX1steGlUg6T8GUrh7X3gHPESt0dd
vcFdxE8yREWH1gjriae4YGfKsKm30wSU8KJULjNy70hkqPMkFGQ+eYuckHPuhAg8kwiTu4yWsTi9
wM3pJM4+bUIJNTjhSSA2L8+dssa+SrZfJ3LwbwA3UTprpvwEfGbyebvB5qxxADeM01DCnAFMr5Zb
u8ve08pV2dlSyCaszVnUiR0iK90iVfPZKcpwfwoynk5pFJau2O6pNUi7EaWO/srMY86Z5iSygbq/
jSyQx2GpFfVX5Z030Uy+RAoeAe0pVC/QkBCiCL8OODgNh4gQPOHMOUchg5Vl/rSjg/vGm/sPCHsW
l5ay982erxoqtWrSzYUzic1+gNcqi/DhFMXSAf8Vhfhm55Os63p9myiWftjeg2zxqIZ8kEmgqRvq
CgG6n/v+JVV7vkH2SkqnZcHP+7mPOR8XcAbg+3J6u0olGbhE8eRSzShdzpSAPde5LVzHHcfH8ZlJ
naFgTXs/zn3l4st4UXvBUwSfXXgYmxzG+AUsUm/gnuFbE0oVF/7aZQ711uF/VNK6I1jGPM3rWzqs
MZt6ZOu6rqD8xQvfoA78WbOazTWrNaF8jqSOBpJIEuo1LR3W0Fms/miJPCX9QvnqLEI6+Fy0FJdh
bfXkqzNXo77V/AlO23tE5gEEse4hRL6u3riYIuBruoHad1ar7Ot0s1f04qrpDQcI10QL19Q3iaDW
T38EnzrjnFBPO0NAdIOdYL1wI5Uy0sB+ntBcx4JF1nGRUiAhBeTKRVhQDE+v2yFYLU+TJb8K2Wyp
YgvvdRhAo6JGzeV07mJA06zIynOTXcDs+ZvaYADv9AKrADttyNoytIoxZ3lFUPEq+/C2ZM0QBydO
9Dk6zJiAR1V865jv9pcXeV3Sw8HHIsZ3RB0QowlspFHbXqPcNJEPLrvyokKELbo9cXgsDfMwIgju
Nq3Itx/Qfnyt5dUP28vgLVBtOLuNDivWN14JHHiyteNxfzz1KVlpClmrbCFcK8MtnUGzgY61H8lM
ri0avgA72By0fvMHfvwUdhu/cxTbKoqbSL/l7og2x7MG2WNmE+/EZlIb6FM+RRGR07+I922tP+0h
uvr4onC+Gd0+3vQ3iMg1L0ZxY54jwJd46F1KkLud5KGQOXbxWi/LHgKiMXTBP9PNNkHddeOZGvlg
4PcVckwqS080E/nuZaU203LSHI2g/50/B1LDnO05z6d+XUrQAd02CBrIPDfHlLjvt/cJpOxz7h2l
o7VhAJQnMIThe76wMcRHKbDczya5snSVedLmZQAawQILTxyzbtVY1Lj7debYtK9Q9ZQ8sx3YA+iV
iIBsvhnstUjNk+SltSq2xtnEX7W6uVPMd68pZKX2wnAit01hZM35oOypYBO5I8pqVTa3BvbrNhAV
sz+Q93a45+9tTZ+dODyf+8odEhOrEXDDdh/RNnHMda2WQfRdsMH+jcbMbbZ+5T8bMOlXmspBwyOH
SF7HXmG9Qo8J/3EI1yf6GjNZ2epuzQLx/cGPrEw9LgrsWgxwWZhyi+SY1ZjGlouPRSuOpnpq4MF7
snbCwsZJccwlmQCWB+wM1dRb6o+NGU+Z3ySAp9/d4lvXMKFNIAJSI4nQQ3e+p+Gw7vrDskCQEQEX
3e0Mzw0++jPwuL3Ql9o460zdgXgnt5p/vJzOxfCMj0+5XvWVxijEnOTtGgq+Li0eCwub/ia95d8Z
eT1KZoWo67d7v8b5tggWLHOz/W/dNG3D5+Opt7aGmKtid7P0WWnK9OHlaN/Bz7FF7SMqaPvHnNgZ
g3Y4s5PIW5NATBXaTTrQ+O+jnL/MN2ld8MVIOmCvh5pnfeNcj8nT/lDyh+mSDxnuW5C8iuB+QCUL
RRWEtkz9Qc7/+PlYrkjjD1fw5Rma4SM1KfmEj8Awpr+0G3raD8LnZJNzOPyPMfMpHHE93Ba3D2Bd
H3yYE26Cb47eHdRBQ/BpHKBP5VD+FfKMeviWhwDCr8hIA+W73MZ7OQUbYxqGyhls1luBfcbFGqm+
zyiPRCCiFOZQB31DqxBFNHEfMsFqUVdIn5qm1MOjz8ksQXlWvRAgt8+ZaVSavApf6swfG82kyzL4
jJDPQ5o+ZNomX5SFDw3Y4JLoifP4VEqzNGlvbxtajISFu4yRz3wePuz8g3Ig2jymkDLxSiASJZe8
4D8b88F3cUh7wh8iH8mVVOVlZCu53BYVrskoQfaXkICdc8NUF65i70x1H4AShaqsVzk1Bb2I+/pQ
NpiYKCqXrJORBuGnHAbbDoxinG0aDDAd5ZKunHWpfJTNmf/Y4SHmk0x0kHPTvWME3FJQBWFUdBI2
7QRO7K9nI8/DrjJU9ZC+mdOal8DLRZ1jaD+jQ4ZWLH3kVWmbkHRkw7KqNcA89mrhQWvj7+EN9OlW
TfWCGQZV6rJAnoU3m5vL0NDtKd/+9kUQGaYSOzmO6EcofSWm7woeSJGiVVrdUuiVzSm7yUEXmPOY
iw7/7+vCoW81qvBJzggUvW5k9y4s7Brx9t/alPw3cSE9aKkDa9NFSPC8+1lT8MqHdJMYn01qOlPu
RxcH1WrCYBdWRUcAIDRScL2ENNpJlExtQbMAsyh+aY66ETI4Cn2ioeDIUmZ3tf1EoEIEol+u0qGC
HSc1khrTHXdBqNRlGJYMWzf5mma6EDiw9BVhqTWCF0JYEW/mkK7Gh/WBhKFnu95nUPZRRIAW5GfN
JiqUPRwQ9nWgWOucAmFdPMjRI4UHp9SwyUNhpD6ssuNmm3Upvss3jLW6/a1GzHxjxE+jv6TDv/hD
//oi8SKkMtJ3Yrbos8FJaHxwu2EpoHzoRCu9pWcKzcCyMANpgDBbCgSQvRXUQridM85zC/X4XlaI
Xz1dXuoGOHIKsyMb48hufjyQ+rwCIK2st2ha+cje0K39/KCflTZBfIXNhkBb7bLfZDlP1a/vli7g
hEEjE2CwbE9Mu6WrLMIgsHG6tYOo/dxS/NtqdI6DlJEp6aVO9Eo0KWfeQpt8Lw+YQpmwtgUpItJv
1ncXyfqZCcDSSaVzIDax47HSUj0j7Cn3g/S8ba8qr0fHMIiwNGEatWsHqwRQ+/e7nspMdHegCQTI
LAPmTctffx4xOfbXibTGCtVQuaXkxjFDsAuEHYp+F25WsrPRDragFyyjg0S0bjS28SdF5nDXohDy
zxUrj+0+LtQjg/8gghXJOswmEysqK2SgsFBdw/oFOncnnfhfwp0ZBg3iElB7TRarR6tuX3IY58gx
qpn6j5bXsNtWfG8nUQudvKKo//Sp7bFrYTD6tb1c2FKE5cSr0Y0VKjn34XMwN7qy1zuJAK+6aXJT
1lV/DKK+72tR/PoTcmn2SilojTuvpQRCIBMQShi/QkGoTiaCEV5/dIpD1asfcsCK8NarEuUQh8nz
nuN655/VDnrEMs8GcasukbT3LC5ewIyelRUvsT6foH7S5X2Ng7Jo0Zgsg4UYdNi/BkvqEjP+oCpq
CItQltpekjA18RpEqKMrT2JJSxW70kM0/8xGCpW46Odn+C7wpVfDm3cUImL3AF5gQd+M6N/+a/y5
HWupIiE7mBk53B2ASGkvk635k40q7ch5fgqEbvZQT3M+Ppk5tJbugB0BqCu8maGnHDP2lXPL2WGi
JVD0pbUgOUOiPNBSqnzSUjkOx+irnOoNDgpXEFll6xRaYi44zq8zvi049Dr9uuYLbTQ3UabTe9R4
Uipbb4QdomfIs+L0K7ENwO/GAq3+/OJ7Uh0Cku0mvNEAxBrze9pc7W5SBQDuXWSQhzwIsNuEjt5c
0DSv1VzvmG1DpLohsa2LUCrXZLVAFq0M7DMtyAIaHy0xWvFSzm4GoqPc2quKPEuanst/Zc5n6KwR
5qrXlaoxabeFRWsp+wvq6RqAyfhjKmT4/5kHTCrHhI4EKyZaP3c+vavhjCeGOCNuUDILI0iYNAlu
KX2cNAvV9uZE/ubq6oD/UPCHn/Ps4z5oKBnUm+ING4S6vAhTx4tMrsV5YTON11wICnXPsmWWJTiw
7xmtDNFFARgUkuCCMTZzhieHsQmuEgP5XR85Agl+GUnb0jKCXPL4rnZ+JYeRFK/Zu5WolQKq2Yqq
K8AyILH5WLGYOkF4Lwrl43EmuG7PBpaLHajopsvXZBHyD2u95nn4ahdCR8YkIscRQGPbtKgu3Iv5
LRUfJnx32kb+cWWGu/znwu9xdZMLJ+eKZnlw0UwubSFyIhjgaU2YPRFG/+B15GRmm830SO97RBQ4
BwNq/+r2kIFUGnRHIrnlo4ZEYXgIK0trmHvd7BbHgyzEgFH6poe55vgOf6hqH0AmwfUqjpFcxX1P
S4HsS62a/E17AYvb/L3wTyUjm+M79JhrTjCV9TFnfr0au7stkMaLxiE/GTj9kyxnhLp7fXMiN0YZ
wS+IfK42AG7GrYdG/6FK1DNU87sRRKdWdmYtstFN4uB4mn/AXgeHDg2FVgutSjw6iSaWPOqFj6d2
2s8O8U0Cs2FTwW7QccAU55FSqBu1U8gZaMmzj537fjzFshMzuzC9U5+/rFbifj5F+Ov0d8hs+Eru
787WWK+uvMecsTKf6D+8n4r3Mfqq9ss9gjwAuY4dPbOvR4NcZ0HQUCb8xfQhqA6OfZoOKyyTngDR
VDUrLBBEe1l+JnUcwNwk/U140X41aUcwzrFyhffwXLiF9Uzts5HE5ij30L2O95oYt/Tm+EEw+7M/
seoaZgbiXiwLsDmT9hRG7xUSqM3NH6ftMcmUAYuRHgGb6RtEm2FKSJ6Ej+yy055t+Sx2ikSihUvZ
PWAVd8tkEYC+i4/qUjzR+Cs0pC5QQiJh73UAAr/d/y+W0Uo8e8AxI74bTKsTSclXtcB5WoZCHQFB
ymgL3J9kzssnsJNEXJVU7DLzxOyGIBbQPWxyPUZM0nLG8LF8OJp4t4rnxfSE4s6LddGvbumC4eFp
UVPpJtHPRR9E4ohmpeGmfQ2gsFt9OfbPZl45YFTC7gdMMzGNeeSTVMvwBScsmapIvqjnvYpowPJN
/KmvVsFLiwLMvL34XXgBLr4svCEHhOIUv2CPx8iiZg/dG65myyzRRmjQjCtcQ+gMEPm+791W9UQd
b9LDjcp0UEQ+O2JFeQ5rUFMOhsxfJNvbZv5r45IEKlGuaM07lgBot39Xs5qZwDjkGFaEjr5BB9c8
Noy7NnP5PN8V3u/xl68ghOnrv+FSUPdVk7wD+W0lSBkhVtfTWSbG9dQXcZctDYMXUdjGh0AkYPKf
tV1KYOfIbNfnIk0N2+Wv8Lt28k5yhlGmPrmnW1ANf5BwaY6hqDdNy5XPwrwc4tKwP10x0SW6JGZ6
o6dre7xJebXbJtxSyiKjt1fdVQQ/gcOQ4QQ6OXhFex/4laW9DY+rwuEfoJeSNQ8jZHC2fPo11KLq
1cDKUnV+yzreLJ7lfzT+TWnBjfDajHKauDsT0Tryx3S042wgb2e9QFd+JNXBEg8Zn8IQ8r5Z1xnF
2/qTPAb2RF3ojTGTgh4oA6vJ+onVHnzYY/+WYUaFEMYo04puzQkFRaE67j83FxowMLgebySgja/r
qjGNpdq57urto3H1ZFENrkXgpSXww3YBKiTTjJyyuWngd85ubmhncs6nQRv7JekdZ/+m4gEZ+eKg
pFGgfrxTzqU69PDGmI9lhRfXMMpIt+Y5LUt8nM4GeEMWpNSKnzRKX/KnwtPjg5HJit2A7mW7d1pV
nDcYhJ/fKi7zclS4WUTewd3hE9XEqRLXz7ReYdWde2vRlYwQ/+oTpwdq31g+aNT/jcRtPw998sBo
dXKfHCymyS+OtZF7hEdRy/tvsZeJ9/hwzlOJvzD94wStr4Xx29gCmMMnMdIz/btzhxBeaDyTuscZ
TiZ3loQ7ysYw2SfAESu6PmOSZ/bopz7LOUxP1IOdnDFETARCx+DVTPUQ0ZIq9T3BOwMV0UMtqogB
RYW2OdJqzGsrlX2wuwZksmyaHDf4KYSlQ0HLFjlWDqUSWedgOeWcSjWPz5UW+dQW+g/VPYTxqTxp
xbRKizlmnmM95g0QkXMY9CTmQv2zgVK5xj+p1ewUFnyfFqbPn0zwfRi4HBJ8pmdY8ficrDlFFcTY
vWXYB/or5g2f9dGCJC8S/U3CUQCY3PCuFM8O/qpWjF7tVD/ZLHTnl233SqybhpL5fN7Iwj8HuSpe
NvU9PXNjpnTqNUY7pAtR4L+3JC7PqUYvb2c0ePm2RUN81kqOcdk2LQozt9hBJYZuF1mJZj1/WIo0
Qi7GexYPDaAZFIgDFZTihRl530mZ1LK4q6OCQ/9vmFybfhGJ1AQz6RPO8kVbLnPYgvj5PbFMRyuC
YV5rrgbbxFJOA1CxN3MiFMh/oD9qh9kjmck29kPT6kdTqP58SMrn3b4jHazhuL1uVW3TGa2FY1H0
dYtEQHb0yxvY1oyPY7Ck5h7Blvblty0i83jj9Wr4iEawWBuQ4eDGKLuGPSW1Ggi0at0DtwbekDWW
4pkHonXMCVcmDv4lTbmWIS4Lg38wCGE3rF2BYP11pTnnpVUKAkMPDXOzoVwQtEDlTmrEGDleafh2
FBzBQsXOSsbUjNZY/8gqVSL5TW63gZiwslECscnMoH+LMIRuu9LHCHvHHBbFqMBTpjyFaE71SiBx
jHugzRh9qN8JKE58BiWkcZFMZMV+UOqpZuNzOJ0kXUxRjvxM/pX+hBjtK/MLeEDmsHmGV55hBnFa
vMeF0v7+hfSZV8H12elaSlVvSHuMyPWPks0xrF3cqQWxVVOW2HnInAiD3pfae86Yco+wH+su3szS
Z3bNnPCSEfo58OW25T7zLSVXcg3m1IWSjEkFRTM8gAQGQ95zzB61YSlQcQZW1H7V7SnEBUOpKaql
IzNmiZ9rd5aeJ+nNMc/3V4zLdUFhiDGW4jGn+58r3VrLnmK6XmwGrapv8xtRXTN9bJEnwetnkPfa
gpArMIuIZa0ffOu6GbV14oADB/qWf5b5osx5KA/1TshT/MnC2Og0ZqW4sRBvH2qFOQd/HSOf4ojy
UHErn0VERI+zHUPUJC6Z5mtza4++Yl7o8QdBdtvkweyAll6hFjlNF80CLYWd7NU95TR1w3KOHeP1
VFVctstRnFzGcI1OAc+hMscrglOiz14Gue3ekF5lo6iAOy7aeHrlm4/NVdvU4MorznS06tudcaAG
fuolyxu8UXbe4QGdM5xTxCQdZhfJzqZv6EGMBMhx0qY0CFC9LZvyLwpNLRSGrNsdcCP092F6SfGh
Vq0dX66IXLdS4Y/FUxQ/V1VYwxvzfq6sF8p48a/TCvrKsnH1/5AW1EKGOd4wJ2P4Po4GD+bLkVr3
MBQ2gA0ve7R8wm3s8efdcwL5hCnvlXtB9q2I7/vvzGvAl+ynGUvkIY7w014n8WELCb/vRaAz/juN
DHdkOlYrVCF4o8ZE3hSnUfb06O6GFn9v/WN+lreEhcAovChoVW1nayT5YJ7RuPj9VcQcHQXAqNEi
IfHEqtUdb1+pYBLvkI0lgQCPpYXOl/7CRR6cSH9pMNLq+hpMqSvvaNwfr7+PGDrekO6rNm3ycvfD
p76LkVgDEcaBW+j49y+mWWAG+9/qvnA6QdBr04dECIFNJRfQU+T01vBO1v4bAeuWTl/4g1odorg7
T31FUEXj31/X9m/EWEC9EIXdNrtsTzBKeJ9rQbQtni0kAhdV/zZ9tLqOKR3xup3UBHSBQWs/L8ql
CyIKPBFK709O20YJxhAgvNoiIm+l7nzCQLYWlPIWCMdt6NO/kI/9AjoLRAqopt9dPk1gxua/QOO3
QzDj9PhbnBfXE8bBdaSK9YUM88j5h/8b4VR0jeTsLklU48Nay0zGq3y+8J7qmgBTx1rRnlCt36ed
CSrv1L/TZOvOzfkkNmUtvJflgE/SOgdVrhas95p6XmSdR/X3NzQOSS0BLEEE7LnYIDwSYXDgf7H7
HOzkCovgBA8QLE9yyjp8Qz56ImKX1NNi+70SyEXXLVhp1CTsK27ohbbW/GHZ3IVaII7Z4ov19Z6f
SG46iFSjKsq5vxFpWhAGUlomuo8tVY6mmpQvzu/XWdE07W3yfnQGtzIXj9eMBekvqzTcW4vpGE6O
DVHNACKHWRwrBU+WL90PUKa01yVvY6ngbWKngFR+bhOztMdXL5fSgu17GPqCk87dj6hWiokxZ5SR
z/ep7Waus44RxkZoUl/UCYAdavQABTlTVE09zTDZ79r7izTfoO/IRqgF5SbuqPVTw/8oyPjI7Txe
PVvxDoLHd5OW3rMiAfEm5yWueAHui36XKEL/QM4xU6+R8uupbynFEWNuMFYb1dg0ajMpdcYGVfOJ
8oJmb/pGCTScD7zzscdDAt7jEdRiqRxr6SF7c8i6TF46NXnO35sO0AiHSv3Yd+vd9+M9tyrvllF+
Bdl785b4Fkcj3AvyAvDlCDHfkaykAAffqrGIPBk9Nz1MkT2iZa6YwDX2Zxg8lB5YLmj1fMgV2SxR
/auK0sCBc/pS/WfIDmw9D3dSV2OO5MMW9+p10FuOwugmpkFbtZ+OMqVCUnwz43kxVx2pCXs7sbhu
PnwUQq4kASJpL2IWzEpE2CZ6tmgjgu1n5A6V96/7M+qf1qNXfuJ23S4glJdVa2w++SvseR61FlYl
MU4v5Ggww/vKT7aHi2mBFAwj6IcOzLGAuZFjZ8+C7Rpxpkpnw5E0o19ybiq+t1z45P1FQXV5Ugn4
Y13Q6uA0u0pWARR3bW1KwFFhRX84vB26oSISszcivIm3kpdFlc+mo+igtOnMXEBvXNM+dM/7GTOS
Iu4VacOGqtX7FZ/W8fStKHy5u5JvvX5dgXBhAM7D1/GwzJZZgzdoty2Plov8+op/2na9f09SLovj
vi/hfl3fV8bdCXUuUK79U+a+MsgpJCIYdd0YaWpLkye9ERAzJ0/s0E44Wo9mw5iXK66vkrFhktGc
v1bAsWLs+g2cQb88YAxa1jrFMmDfhBqbgZ/2IWqzMFSvQe5niLLYFpsNKPycgQPOqRii16bqstFx
h3sqO4ByTH7bAvVuclF9rk3LZeLtjY48I9dP9jBism6VfVMi1J6EAzmTYO0PRcvSjJMvIdp29l7m
RDkFzKh7RUJDk/JKgNOf6Hi4norAerK7NlShl/jPmV5d4FQjAFHygKnGoNTZeY/rofX22ka8XyBk
WGOLI94j0rFgNDd8F1FWZxeRMn5n5NNKIX8sAH6niciuAU5INkmK9ky6emRkwV9BxcHU3r3Xo8pi
nC+tWanPP/Y4RNnAJCPVd5HPKx/6qXFnw7JQhsrQINiJbLmQrgwp3YcvEsr8C84YhORepk0Dje7P
1ZpKPt3qW6gc/dAtG1uUm2YLvtvyIAS/y6yt30Rgu8Aa9hZjMtWkVced5faUtsdYOFxcJ9GYmIgE
k1KhSm3KRnPafA0T7TCqc2kqjFQtWj8Ruyxsq/Fa81rOuNuXia8pHFRzyO82CIb1MzZPIm/eWY9W
0jvHBffU9f977C42fEBZ5MpC5ApZs9iur+KB3ecY2NA1i6FCuOek4XnxFyy2Wkx0k2K5ZhigkrsE
VRuNHHuvxJJs+x2eSAEcrZiGAFNXgPdlISAwrK4Mzmh2sBZSBTxGirde9lZ/8puzW0fnXdzdSNB5
CBVG5O1aKhJAAxJADTGfyme96vlPKPXmG7DCPujiyUnIGusYMQL+70uGwhasNVFVIsIe9HQGRrd2
YBf+lENX8HM0b4CsU1xBXIRdjVZIEAy06yQe92LpRia9CLgfVgHo/SfBXO5+N615v558pXOhgLJd
tbrYevOrLabOO+1tzkNUtO9FBOkGERVW2ISyQ2eAoex1YSttx8fkWCAxPWwCDwYUkA/YXlv3iwX/
Vk4ynRjecp8U6ZwXAxyCZSb8cZQOsqXC/+uT7RoU8+pSu9g2AXrQfKtI/+5JEiK2RFfEL408Miwg
Hszf7iqVtTXBiXenriRB4GY2A16AlJhuTiCq14S7wtZlpDLW3+xRoiS1fJoJI5BXE7PnyZnzOl8n
gIWL32mWav/Fb6474Bg5FdSKIK12Fw/6hpJV0ALsDQ06lHAlbmmXhmEFlzBQwp+pAKCTIlbrRzfQ
KKkuP+9CGSzbv2TeAgdiq4zKrhcEF3r4CsW1cFoQBYFP/FjNuLTVcNAkCHz4a1M3l94w4JnyQOCa
hXvzlykpgU7GXdxlHbBMXSrNGHTvqUYT6BkBiOrXfuEymCbC53Flw1+SJhA0tZDmRKA78vIMXU8T
iepwlNiOMEaN59dshUUEbeyRYUj0P2QfrSbM4Rj3zCg/dWr49nPwZP/pVUyqIF+9/BW1wYrrOUzK
J0qNlY3jDQSg7hYspKrijeuIY92cqdGgRHPaEXBKi1byby4oWHCepAUXDd6T0aSKzUqxmb3vgGsc
xiIJa9WKQEbxBVtUGHUt4Ibwu+PIKU925rg1ufnhYWhxxpGyQUiovpLs2ikVQOyCS8vbgAf0Mls0
SMgZmmAp+x2y+hQ1kb7GQG/JZOQzmjOTlvLUVUyKkkHiSagRwBJVkv5GVJWyWUu313uzSoWA6ofo
LQdsO9+gFxFVyOhZD5hnUFVYS/8jLI883fL3Cn2ISI3DGQ3coFZqLx3r7nfjyuoLRY45oHgyRGbo
4tQHKZvqRBUfycw9rXyTnOgEuf1ynHtORGuyGDODWe6LWZRQcqydiG/BxOX4TlFR+yXwMzGTb+Sn
oUXTXmwfqmKpTwEoKlINV2+2sWzsykiCZoAz8iSJ8bZ3fFmEn6er4E2Q21ubCXWg2VIEnkLdf4Kj
XyXZyPCPbApLzOsGqQaa0G7PCmdxL/YmpSp2AfL51Que35z7YJifhXXKYHvM5qulWfU8m37LMoL/
RHtJUZdwMDY0iEs7V6OmwPjjJkGtgjP1w+7WIlieSBMCa0HYUGPmgDxZhIIL2XHjwZM1MFzq7cPg
4eHL7lh0rzykuTrAWQvzMc8PJ0XIw6Ai25ryovA9GsdxWpYZcIUKdYeReXbhKhs73s25AGvAQ86i
flJqKSx4N8rAIFYpR8pTbOOQT/ew8Nh6vEfPFaH4c11oGSi0wpsp/lAxecyJkf2UIoiuZEh1weC+
NofCl5tMXhXisa4hIThfUO9zzHEslsw/HBEkwrNXdYYLeWLM85I58lkkvz5Ok1PL+HaGe+Il7J6Y
0Rv1MuRKerhZUXqiYStY0egwoKG2u3AYiH2VfG6Dp6F45c8f3zUAhasX1eszSH9YdcJhYX5q4rF0
HQ4ZLDYrM65zYwXlmCcL4YrMEMt+k+6qspuXt9kgCpu1PI82KN+MEOPrYOWbO6OLsy1ef5j+RCjA
n1PaHCI/+C49q0DW5T8af3RgWAuWDCzBf/W8lpXIq1kilo8AunTiAK+pEYGzW8hR9NouZuuQZ+A2
nPhiPhMhXQDWqg86hI9f0XjxtKf1UP8eDgyScWLJ6rMwDAhaVo/BGNRLTx4kB6jxOW9l9/yOGZcA
2lUUFuFKKe99PO35vCVfGqsq2GEPDNH8CgnHzLoEsye+n/PE/i6ukMxpl7SxpeF0HIDUYPnzmBO2
1MqAK2YBx8+aPZIeoqA0avBHPn2Lv1Ig0WHy8pbe321FsKJYh2nFaZeH4+AhiwDgp4JVg2YtvPxS
1OFxB1wdCWIL/OJvfrTy0/xK7UQ14is/Q/dqs3PRg0/DlEi07BZkkgi1GzE9SZgyRuR4woPOMtcg
Fiv8RSh8lMHg3tlWqoWE+toJ6yAlz59WM9+t8FncUJQjzslD0ZJVfB3LBp6rAq2MRXvGjQ+y4ipz
SOBACcX0QiMIv9FlnW/OCSkUrNOOi1hGURsf+n8uVCBGkCa9OjeHK5a1+VeROn1EdwIYBMAQzNRI
dQArfaADAu7qrtRuGJ+AlYpX/Sh8Lht+pOgArczj3xvywy7Rdoz7b5LSc9zfX98+feUaSl6CQJ5t
7MYp4Va9DSkKHD76xSee9hCuG2bmiQ/YhloBSeqy2T0frbj9E9yK4562Ssq9shFad+jSVI8+IIWt
XOIrRL1KKTkA4+xmCgtk1qaGqNRi+UP7tcyKDnoSfUhonErWioW7rWDwYdgOVeSzz59Ny/hE5aE+
Zpj6LA5fUrq/GJl/YDmVEmZvUK28oswzWeNBe8SWEJs2A65ccgYkAnw5MOgfV5abNK5AZNWijrYt
2GMW0WADKJ2C6zE0/HenJGuSqJFTFbsw03LK66op4XhbQlzeAAM7+HjkvZK2QXTenncOHT0poFy8
uuGIjvmqA7G9SjgckPUSYPMNL9jyihrtgquMSTrVY8SBpHXHnyIRMBvxt+nehzZCAoxmcNeFcQXB
DTTveuLbaEd3RcIGgMLuODKlsPh6jQXkJamX9yHRKinfNuOrV4U7FAnP83fYDLXwBCdaPWuiHNIL
8ObIbQ2aZpKZ116kGdNvGo+FZ1DJrXE8V5QIKQGnPEJ4yr1yPI63aDfOvB3VUjoTmOvSBNMuvHJz
YBxyMhvvUcIVd47r10uRDUaXDXP2G6R8cJ4hkR6I7/nx0kEzLIjClPvrgmrHhvsUZv6iqyH+aczs
L53BYjVwm+aKYoi8cjMMlFu7JJIWOX8sKk0U88xupoYCvv6q7RSQZQKFLWIONVEtEqWMksrRKipN
JvBOcDxLTfIBnaW59NiG+NdJENUdeRbaS2Fr7vChHrDGPddJ/08Zf4JjC78dljlWqjhHRCx818cy
jJgIJ8sMYu+p+Oxpwi6oQVp1cyQPMiiSMtfvvnzllu8hxjlyTbO9Vm7XAPBfvoTnNTQJh85jsgmu
p+w56DNgFMzFF8JVko2aIVv2LmcbxsAA4F0udJ/6ncm/lC3IjG3iSttJKcbUQ8x9/kk2vsaCnXpN
L16aeA/ID/xgBMpqQNUUnY1XqOsrS2QoufqPeEg6YZlxF+0OFSE6iJqdNobeaxcfvSbUJRF0ybx2
/Nzbi7nQ6jWm47Nh7JhwYAf+IH7brC7bVspPUuRE+svdgiZKxl8W/W3lgqnAl76txC3w+SiTx22p
6ka5h48wOD4Ee6wCNuJV7GhG3ywkRUhEpQLyrkN/IbpuhzwCEwlUa6gFuzs6uEVLbQ3fnDHjsXqe
J/qpsJHik7qeBlrzOVDf15VvbLjtv+OIyhlaFlPpdzVg6AzPhIh/5R/3699xl60yDhArgB2IXmmE
0llELjKSsq7oLOXYnjj+PlSMFc8ppkgSqOZU1M0HV8gsyy5uBLxGVSic0R1KzgzD9mT4qhpaM5Kh
pTZh/12qtSN3uiz/NK+TcrvOADBu3gExvSXJI+//qx3FCuHitzo2SBMJPYjzEsqSFE7izFMsbjKx
0GJN98QAwclk0Oy8vpbTdmG1psZ1R48/xUqoz75k+KuxW2EtmXyN3CZYQWKtnusqFqB8nM57SGAb
e07EZxATZHq60WgpILTZRJHFaReDsUZaHIWx6UaCQdfU/fMflLj/FcWu5VfMO33mRX0CDOL8GIMB
Bqd1VGkZBL8C3u9m7xf458L0VG9VeazA2yTUkbN+IOU4tkoWOAe46MwSBdiYqcZgfb9y4WzspMLA
rd59EHqIB/q8983+0EyY2NJFGQleER4QF6IRGqQTdOZ4yorVlLLzRJlFHDyK5tmD8BqK7JC5AIyX
2JQ4ZgOnWfJ0oId0exi63LohirknoJ7wkaOmniy7kdywKxDc5u9EFm83YFpSZnoTI7SIYgBM2m13
5SPFd8DcDFycnfGRG/lIUmfWyLV23W1i+QH9YGTYw6X+iCRmORJPDh5YfyzMQWBdjJNtEYSKjOSf
mnAyq2v2ekF+R6K0DvH6L1nXc29tlEPqU4za2rPa7Txh2itku9+aNWP/t+3WEwsFUzQoAgxz8Ay5
wPtpDJpsX8zJHIqlnbOMAmuariNUSGMjH6+To+X3V4OVWut8JdP5ZKwWBWOazwXDTd+lq9HMSYTb
+gHnHWMh2E6IlfBzMfAV2JlhGcyyJgAdD+rS/dywit/XQ2iEfYdp0sKkqmzo+qGuHkI4WA1HtjKR
r/YbSaN28Q2J8lKEPFiz2TtICAg8atbgR5rxUD9Gr/X2zFBGsr6k5PRhPXEL4fYb/Su2A7diXuEL
zBsyzHmihwTgMpg/nuVLvAaOHElbV2utOT4o0IpUCJe8ueQKIdzjyTb7vpeCHHxMYYccENXtBqb7
nbnpnu+2EN9TCFZmnNek0LUIn6wbcZMyP3GtopdMpLY0kunKsgCyNdAot0/D9aI8llMJXYSjD8Xz
EetImXv7b/S/6CTCjLg0wLScsFRfzyi9u0BMffvWjwlAm4ktMgIF4vu7TzTSUwHSlBf31LOrQK3R
pM5fGP2Xpg0xTLdYboex720R/j0QR7Rzu0XAxKuKKe6edL0WLHnMxPl7V8aedf3adgJKhJWAgDA2
E2+rggLRm881jQ899olDFnwe8CLDbPb5e8M6CeSQtET85x+fqoDgozKsXh6fOJPnz5v7A34flJC2
PCDIgo/n8MDXdpxxwFgJ0cBScSczbfIwYOZpjEt9XE1DnLv+b6tg7yDOQJymuruHcK+uCnIpu83H
adKQM97h1NMSMqUAzVxnZvzFz6OImN2c86LdrLT5tEihaDi7XfuJbPgE3wsrsh2EUyrak2YMegxK
OzVJyu2DknB8jb1F2b9f4qJeElqlQpV7VgnyVhYulozlevP320VO9pjKtDFWJ105W2/HWo+FJBr6
ieOmEYxtzo6XeKf7OjcbXGojZzGPemc+WyTZmSuQZzItbhLSEyWUn5d+9d2zHq5icRZguprBnq7T
u4AxkTTZjlmtmATiCsgAkG6WVWxv54M0id1u28LQsawnF35bx92JXxc+rUpJNZ/kG9F6Pe7Jy0MU
tj2FWLq9h+HdT6ZjNB2FdYyBes4cF3U/JvxploCVUItTq/IecGjtWhQtcoE8EXjhH4vDcK5k/Xp6
QjC+W/A2nxxwg8vpHl0Wkh7mf6O1C6G0m92773v+JQOaWGX6H+K3LXeB5D2Qt3jk5aucjVzgk3YM
PunZUEkhm6g0lUIgpNYV8FqewA1nZbxO14c0yjYxjbhVeuuT5L82XoC5kzoVCrmCQSaAVpmDqTVD
++ekBA7gDWnOnLkEM4SUJ9fkJQWGtx/Fz/8oRSiktnPRUQuEnmLpS50K9syfslUzIAObENl5A5he
V6CqD3UyA2pa8iJluyHxv26eXsy6I9+4qRsfbr1V5RFyOY7qni7MCKJaHdq/VtMbuyTegFMHSm4y
OlgwfIEIuSuE9oWpMgT8oBp62W7JGWBEYdur9wOeACyqdyccENXEEqRUqgog33goHtJTWff38fJn
sWsIDyVNwYH8RxG38iEPJPVvThKH2Wj24FzDD7j9JbDaSfWSxauOBdsgIm/S4hzxyT0a+QMo3ziv
ElSkGRmuB2T+pxfJAQsXazUqV00/Ojs4f7ZuGAoWRLVCcPbs1DAIgnMKV4p5qPMxjO+m7HsFRJfi
DYwv/5YNTS40fnClEiFH8Wo/PQiKg5gNLOwfBB9AeFT+bjXTexOC8T6UZmTVsKGUDMf4xmokgkPL
HPVJIsYPt062tz+PW4XC4l6+JTRYN3zrgd8egMdveGEm4GwEP+ruuAeVR++QOWdHVjFm6OA9+W7l
5FFDPu/TBI8/3Z1rUtjfCpP60HQskCI8lbM5mHOTHKxCb7vpjM9hFf5xIzLhaQztnpdvae4FsrTK
dW6KmmdjA3vIjtapDjyQKUSe2aCHLQ8QLar9NvU9agkLc6zrkprLc9qTETJceyHXdtgkwlOLPE12
q8o0vbifQvSiC65OZQM/pVXA2f7/ruqXrP2Y8mrv9Xy3al0hmONifNgfx7/VgTwZAGBS/cFjtBCs
YK2TxquTgnrFfc/HdNZlYBiAjFccfebLKXEuERh4TgeKCLQAwje1uC7XKjAPo5g/Y7Ov0X1uWtyz
WQYiuHdSVshMGS3bI5vLpdnYY/uciqcGeuCX5SnrVRQ/IZyM7Vc9hXUaBqyANtMdFk1u+3rbD4N7
N1PBH+EaenxMIA+fwN2lwQR+qkeumHueOZJ347DALfMMZZtpJP4FI57OACvArHLxXd9z6ebZo+jX
aGIhL7gJqyvcyevEF4cgFwkj8Dcfo6yufg2JIkDgaZm8Ecd3vr09XXWU9Ubp0+ogG0I5P5AU5oEi
8Cr7WcWlusGzGZJ/YeGrp8J0UG0swuQq8dqKfGfZiJLgkhD5q3jXYPh+Xs9om5t9fHAMqdRVMYnE
wLNMNlP3aRD3/vcVoV5ysxmarBoDFlAnZoaWeaXQA6MAa2dEO9MNqFtW4UwCmRv5afPMQ1TwkgJd
hXXixS0GVneRb3uldnVPriMHml++tk87effXqzvpNpNcBxew8E/F4HRw3sSsCbkzqMJv/2w5k5s7
MqBpg2Wf/GP9xShaVaDrmMkh8FuKw1ZTSKrhWh+BwgETef/fUTWuJmi6Y5PkiEUOsuq8lOPzQSis
UJUCCO3T4TboI5RVKsL6I3QfVtw3uep2cVY3sydQ+QpieL56ipGSoTfNBrxz0pHftNRfMGdo+H1z
tKDWYIw4fQuBIxULN986cZfiJ5Z2UtTzhzSaAJ//+cuaZ9v8kaFh4lYFBLvkp6kSlumojik5Lhuv
8odKceOCy1/9B6rZOyyfsLUOsHGH0p+A/zSPDbZs32BOa6szSbBN3SP1xVYYmmoERREQzv11yTF8
aAyhTWXLAdbq4my9DePxKMPOHuTxpGj6W2m4jDgDkUX3mVqHDdurdSjS63HYqRG1Jd0rB1+I+OoL
fqkJfFS9/xi+D+7AxWdqUmHizdKuFeYXjE+7iZ6flAyMQBy9fP6DFcn7SgEC4VWhh3GXVcPyCKsd
/aj0vTWsmG64+yIjvJV5kZw7Tzt7NAXR50nz27arEojmQI6cHgisLmoOnfRxRW5ePKwi3ZEL5ztZ
sSRe2w/F6HnQjDAuoJLhPTPrYkbiRL+NyfM5dh9LA06KPKdnqsCd3Hm/jDrtsFfL7wFM++zlv1Ig
mf/qAuZjwwykaGkMrwKxyF8r/mXRxwFWDU3YRdCcq2c3odYbPgYPQfPK7OglcPfbO1u/gId9uuXr
RJMxA7ESRjjUiErlbojSIT9hfsmAQl1Sgo0V1xhJ7f0CWPykOu6aM4EvjDTL0jHdDxt3xWRg+M9x
2HcN63i4jaloN6sLAByzb9nKt+in7987GOiswNgkqO3gw+LEr8cLy7Sob9in2Ug7misX4+HPgUTA
yNKYiz2XvRR+gcgf4ko/QXQlP1tQD+1Syh9CTXG+14i8WetIaTJIPJesbPuyT2avVqGmFCyfOXGy
MAR09FIkHW9v2SKt141IB7T/cV/FUXRODdFzAZXaj8a8zcuYE+nu0UobNm9wRy1TFNlcAvzdQwXz
+YRtuFPX2Ke5poPl70E87bmjY722+BzAtHLIXvdMo/XFEUkjfAS7GE3IXpbm7EZAIi3hXMcs0KQl
xr49AaUVg8mbRqcYW7NDh78eWc1fc064wHZDXBjpAfPqOin3U2tYKBRuv/bsjdu4TcDUMT6f2Aiq
OEKDJ1kmxBSBhVAVIZBuMqKiGqZFO2b2beV3/lpXn1N7qzdiEwXRLmThhvq/AarmV14Ijdlfonzh
k3U/+D4GjKo4+6kvw0V6ERbguUQaozCip9jy84mkUT1WSAHp/GUfak3IcQ0iJv7W9BUr+ZNpzw5M
lwvi9BMgPhEy8JBH5Wlyq2038CtUwhvuYCXL8v+lZeqdwjZ4YNgx6xPFzMdZKRVa45gHklAArkX/
8wFom5QZ5va/2qB6U7OGBLZ8XAn5f/tJZN9vzr5bGIFpo/N1024YuXGvVFxokdfqmWjDpxE6hZga
RDTBqblVNd0F8OWxhNMBd40VDrJdTPoou8uRWx9SR/BrWBGzlJTyCiQ/S+8YVZumo3C/7aG9ueaI
RWHkWLJG6Ud0XYaal4w4FzlJuKbTySWkhRMQx+DY0NbAeBpXzthAinzVAQmx5CHcpsSBh2dVwsJR
11Uk62nmBrUdEyeJPs8EmtJzDJJDAk3/vhQdp6bcw3fLoGL9fFjlMLkOJJh4u/Ph/F879duegWEg
LpgYkSo5mvMKOsrt97y+RR3mV2dQ5yNjmEATXucOEQ24DJDIYkSwg8r4KFAOOAIleqFXyH1HaTT5
YvWfotlzuh8LPjENL8O0z74JXM96QMZ7zmeB2eLs+H3iLjNZYI0g9ZsRO318XgLw1vagmAaO5VrU
LwWb9078V9IgBaPY9aj4mHWYyfADVkesKMeA9LxdylzCoIPGMvr+N2BL+lQrXNGTH/oGBfjZ0aA3
eH2Ful1FMHqVGXI4bzOqCoTK5WHjFJmpvvfC90kl/FhVJe8YIhz+Wp9Hgy2V2nOfBGiJJLXAHbXR
CVBFOJUtCwdt04YqToCpt8Bj0dlWN0nvF4afeaDXXfzCE3ZAYQck86eMSkNPwWdPwZ15CJIx2euT
9gbiOjwHrBcRHKqZmAIFF9I0iT69WhVj/OAYvum51+OWGZmSy84tX8Ac3IbD6HWjPpAEPFsPpy5G
JvujgYFo0uWWLwFL5mN9VP0uqpUUIF3c/aYyboCRGtn6LmI5lJtd2A1f8OsiKhNiPl2cMLrq/HAL
ddhUVGRJ32joAChxhPUy6qGQL+N7eoNYwmLSuKLne67kUVlJ18YXjI/uN/nfFwVeW5BAj8+lvp+P
EPrev0b+ya89rVSDq1xTsT+9fmcvnwbrGq1njh8rkIOYBvNw7FCm2bhlcHKq75/BJ83ADKPwWJQD
ascTDIdWqMaW3uGQ0JgtcN2c4FSyaen2wYAwufGjA2cxYeaoeVMRt5HYS5N/lWhuivP8DMOLuHRf
xEONSwPgy8DNOxkRfqb/Vx0etSrdKrdAiO3v9zCg/UPIIsm7L5XeiCwbb22pGOqGAO2LUTnFPHjH
BCZG4Xr6AAgNZNgBhs0LTEXOknCPZ/APXuI3Cdd2NMG1XfBes6uHgTG0TfAQdReB4MM+2lav6Pl5
ObrGj6P5pLZ0P/R1zKruS8ipwUxcOXfi+YJ2rQp+EV9Y127w1GEJqoN/AH8gtqbe3iLhQsCJ/HVg
+nmDdnAQj5ETFjwv719GaCAJ2UT8zb9p8sEVe2P76T69cbARuj2Cmo/e2IgL8W8R61+IN3JHYySS
7iLLk+uQBvKOsiaWtcpgmZq/ZD2D/cCiyUbUJPMIF0/kzVvPkOUmZs1j3Bd7FApGGmZtGz/ljsDs
EY3pCDuRyTYF85FzJmnrrAL64wgBkXtHcWxjPVbJ7GqTH5trGiHD6GWG07MP/LG6DZYO1Q3YiUyf
7GksxMOcjZwFQwfdTSYRzv3klIBbtlsV8m+PHLmMQBLzgpQXf61LwWDLUCECP3trw4kYbeI7U0xU
nCduDUh2eKRBV0XmpgPpgZ/tbftPZ+ab62Vey2IX/eS/havkLPBImydzLeyRsDnpsXHzTvn4k0qB
wZuTs6GrK5obrcw5oaFfX3lKKXD4wiYXhxBDnFXCIDStpzfQMddHN6EYjt6uUxmP1ouOredwnS5k
UGnfzECRcxaF52nXMY2ODTBTkUTzlrfDhGapPUOGPLSiZjmG40qQfLnFme2Dt5lPAPYRrcIKDYzh
hY6ebLd3JWFgW4fclA/EP4gdfgSOIqMfBA9vSsFFAqM2Bt9n9A9KIz8fXZFP14EX5/sbtJXT6l3G
WiHCppV74MWxFbsHG52tUTsLrwPn7VtXyFn5CCvA9XPOC0tivZvIbAyfh5CpsguvJ3NDwEQVPGSi
pOo++WNSuycJdb7p35Y/ipuHueFn05ZqkpmWRXKuv4kkz4SimXZ2W7pXQ3Mnki/IoWlPOtIiZ3FE
Y/gH7JhDaosNmvGymyYl2CuPZzyHmwkO+GpoosmVxvQ1UIRW4smLCfpW0XsQAZDPVMEM6yaW4Aud
Cq2BclkCUA30w0+pIAUO7B9zGZCYqjCETe6/jD26qE3S3fBL3P5cdNPcuKFUSMBw1kP31RIeItDI
0csvm9WNM4CabQTOW5U/jLp2MEkXDm7xefihw7fxNWTjYREwf0CXPPglLlDCRp2s+83xvln3RcP0
ZCW76PR0bijJx5XpVGZV2FekrzZq6w/0+HLn24BEtL4a7opR3omyJ8DvrhZvQLMBc/iu6+M8Y4j8
R1TRFXRchU+EejMIrioWft1UTLPXP0kV5bmzkCZoseIxXRG4sTC5karDwjVfV5Mf9vvB8nSHlwiJ
0Nbnw1Lv4WL45+i0LgkwbMeMj6DXhmHjlTeqcMm88+ZHHMrXJcgciTfPpWLvnl5HU1NFy1EqUZSs
ariLYyw/I6KpLcyPvaeoqyEw/38ynGifrhrNH4Hgvdz8/G7NiORVliNIzKF66/9V0+z7fmsKlQLp
Ef3ESnpwNtYoQHCfZZ0+XX02WPbq/dgnDateXafPxRtj18pCULzG4ARCBl/L1aCJQBeIJBPMHpr4
h1Q2G480NmqC6vpmyTUzxuWPmBhYQ/+OANPoJqiTY9fgXMiTdEHyiJi3ebe/ZQSpnFhdskGER1/W
BJ2JRGzOQ4VH6DwgvXj9VwYxSu6Wb2p51rK8kHmy12Geiwq447cGjsyPyNOE/uUJMDJCPiyCLUCp
5S52OqTpayqXmDZuymTvXSvQvnBzstI0DgDHfDR3ufEhpMr2jXcIVHBC5Jdfb2OTvJ0HXcQpxfk0
4BpBbSwX7Ucr5jcLX4aP8CFj4/AKLoZc8C+HgziuKnBguiqgZW2daHCNHEbZeXgxtGheZ4ev1aNa
rwlB63QoCvXUSY/XMDMEkGM4MMx3oO5V/ILaKyPG0XoM6UlEbum+OqeWcXPqDF7lFKi3JS5G3+fg
cib0OJoKO+deA6w2HnKTqHU1lnFwXJddeOqqZx5hyF1TUT/qlfsOSK+qmdl/l8LYbd1k4zSpGm1I
9SWdJmtE9B4lQ9JwKDNcWQclXc5QXFIopZgefviNpef5BaB916U/UiBrsQuuGB3Oxm5qe774p+40
sr1nu1Dqe2BWgevuotvt7CAEPIfo6fPUJ/kh9lEHvbkY/JngM7gdFgcyObtKpz1RB+0GTfoxqXAt
qVwCz0DlTfiQq4QjCBzBr0By8kq8lzhUjhAkSaWlDc+Fc6MmLKFgUV+TtXPPVfR+7buONVuNTp+r
gf4IjYGjfWjZ+Nj90yn4nZFAV8Q2KcrQgj/1Z1Bs2Yz8ygmZfRycaJP0i/E1TK0ADpekPM4X/1tT
r00G8tZsLgGCX/uwQcayiv8KgTB15/tWBgJKcBEU3DfYlJAJIZPMBq1jyt+E4vmM98cEou9zSQwy
gzesmkkOARBw+LEgbPLPLib4ltqk2jqH1pSNV9H1Reuw7bhRpd3ljef4VftIirZ7c2oGX8jOkmI8
aAM3ZeiWrgFg1Me5H6JtlRmQG/xZqO22hANLihsT1ldEeLdey+tzkB9D8QrHaKeju60OF+Yrtjqk
wgHfPsIcuvGl0en0Cy1ZbTZGeliN6ddCYqndOE4RhalqHsSunQ9He+Lwd1UK4daLFkZjjIPXFT/0
z0uGp3+iVXcB9Pg/iHD3H1OeALhfry6OXNxIVE0SbF6P7KcHv4C7cjXIIzN86gd2KQXfwkTFib+U
I7OBuX2E3zZ1mfkZhTJFeEs2lOjr92x4pQbog8AwemgeDcT3y0uduVaLMcTzXrc6Xc+tKabXzf36
TroAp7vgfxYIMPeIt6qrV4DouOk8Kg5YdgHjI9+UqpIT5bTpqRy9+zWyKT1CnTDaH1LfoRGCFxc9
uXFY7mo1yspmPsOqtGZRAmSBvAZLc9Bd1OYrCVKymE3HXY6TLw8tQpiDTYK6sV5I2wrFi9Dsfbk5
oxW5gHr0AIzhDwzvPeQgPAx6IKzoUxYi1AX4dyjx018k7ZEQu3Btgvh5k6XkieBIlZF+VDvhIHSd
kzB3kK5svuyHnv3P2XmFg1Z57nLK5VDe3ZpBqjbaLpGlrs1YuPROQCRv93z2RbzFNFNYAcbHDATE
1n/O6sAToyWPP987Xysl8jBCjBRK7JyUY+G/gzILfJFZl0wtkFGSMcSLJa9YyTfoKi2CmKmh8zvD
xnxW6cCbOeIVZk8CQeOC+UCXZ0tV+orMUSVi1+06baKrp+qxWkJBVUF1Jkf/h75T/Msc66ENWx3h
lOVuN2xZL8/wYmyKpf4hdeO721WeLa+vBw80DR8ZiwWSXGK4+69EiEpE/HKIFLptjq2qw88cvOq/
rvNcVuFtbtEVHWr6dBaIG5MiK0WJbPuXxpq2nU0DxOZzjiT24b6jiuF0ASUXZbneJj7I7xNI30vr
dAE0p2zmBSPTl0wm0UZSwtS/KNZgbQrEn+Bu2+LnMhGF6eMyRUFmytmI3YgWkEMffv45GWFsW5SC
3PBTDEtDaAOR5j4FIQ6tYcN93yzNaaE+1islRLJMA0QDpNFFtg586+6VV3xPKeSSpoasFdwLHuXk
GjTxgZLyrPm/MVQ3X0y2VYJJhuLh8dM4rfatgJYU471ppBf0/8emd542mILwnSoWacv2F64+fQm7
Qt1PPVoEu/azrhrQy7id+NbPf2+zPcLgIspEZFhLKT+rpQXJRXGXQm0YPuxajpi7/Kf1/V2vC7Ly
mGybQGvgPtdgWZPBMab7GkAdrxE7ZoyhjQqeTTdQ0s19LOOth1Wq41LbSiGRaof34N70UpjF7r9N
/5W/EysKOrjkZBRvKnHVhp7CwglWFJRWb09bKV21CJzR6FZSBupUwdCEps9sO4qlWnY37lOc1LYC
mM/66xeaKknJM5R9R3lW7YjtrmhFop5UhywPmeZeSvcNpcPz4wvpi98f1cJXskXcQhHhA0S1o49n
TgcaBIf1iE49oLAuKGdAJARVOFyPSqWCltag0eBNguAep6gZNWcwPg4ZgwEdacBP8Jym4aQgq1th
wXElyiGE4diuFLLDS2DOvXE9yHwFxVuTQL/FwFxqRP4e0eE059FUgLtjebOUZKo+Vox0Uw293cIs
rZ6kGTjkxm1ADg92zl1LnNDo0t30Balk+fh1zjyPXktOJfp91QomBoB1mLKKGuqa1I2Qp65PkDhA
rLREnovjCpVZSAlCfRQdG7aLCLa0b6ael4Y0bparCGGTCD5AwYNX6rlEvm05UWWsyFEu9elVbeJM
GBGxgfHURhe853c0GHWJlPASis4mA9nPXDrxj9G2AHAAlOHFLMRvblnkLAX24nJh6oDduyJgAHkn
fgRb/Zj+AhWXu40b2g0ma0N1CiaJZbyo0cUqPXpbze+2GEHbK6VsPRtx1nhIh4JsQ4fYNYpveClP
OjKURTxqLK4jzFBgZk5Vh0zEPOzWXLwOOvjwPmm8zR6ZIgTFzNATGiWTCBWsWzOqy4dO0nW6ozqW
ec2zq2QZNqkIH8Xr6qqkbLZLZayJm9jgZf3Whre06xzJ83iv/GQ1PTcXmKe3d9HEr+K8RyFWvulf
NQgmcfwAhRzqdgI9Zr3Gy9WvRCZkHWK4MO+B29m4BSTGyWBPFVS56V0bPSsqfDCAsSF+kDMnIcer
1F1Gen32me5bjPuxXJ9Xhbezg+PsbG7nHyeV0uFzixk8HsWeoWP79CyOS7m7UgOlgeZsOHtrrxkL
+JGimHDrfX3uFLlei5Ae0ad2fAGAQkiA1BFIK1XPKXOYjMEHX1ONLZy2mut0q8TVqe+KSZPbfEj/
r0DdvVtW0s/TAeavHDaHz5h3Ce4eHLYQ7nkPP0dYo2byTgdZsm/Lr7xpzPQmyQSLIqF/50UL/Xyn
6CcMyrfOwvsnc61+6cKsl4trYeTXqWAieSr+4Gnh9njtSdp999MeOhpsbaOMWdrTH82jHEkmSMlC
9fi660JrQiJn/5zeX7/l1WLeLSln1zEBCbZaZO/JiX8LG9FTa0Kq4NW7R6kGXOY1yeB4ST1RSsho
Uc+6UdPaR2IaPf9C0VnEjDiyohd49aJPGHiJsDO+7xX55fXcJQ235HaQoKAKHmzgigDF4oruIH0l
ApFlcsEYMjWyH8h0kMXGZp4gadgZa7y8Q0qd+Cd5xQyB6JljF9GufGK3ltZxjD/Mhm1BMF4f7Dn1
2FSCAImuwZDmH+YSUWbtWCtsmeLTTey6TNkJaON2Hb5iwZ9R5CXMiXX1j/sH/GblfHAD5YD9LG9u
OXB/Ip+YbTYzFL18RzZYYef50mMy1zAsUByAfVc9VLHTmxv/G0rnmPvYQBn/KWNHz3avCvxzTBJ3
I1qA1Pjuq+RI7iYF0So/avT6w0XJgQ90zKexe4jGw8oy6Z6SlX7yrIZwOeE0kewDIoTI1F/je6N7
QFS2Dd1X6HoIx+qn9B3onx3me/xPLrQKKuR9bJ2KOp9SA9UKhRsuqWODWqdy4I/UTCLnUEcGmhho
oHvr1MnQ5AjFpv4nA5BdkijpgSNWuWkI+vAsDT6kYxHad7dz/y6QjDT8l68H2WHpBm0rmBZew1Lw
76E2VFmUu7M2X8ZVnsmH9OWN1kFj3NFThRuBg7C8YX0EWuE+nvTjWaBOTD3o59DS9KvQ22Du3YTU
nuUvGcBzTp3x/up44cfuyLWj62NYSYCEc8sSd/d353ek72ljaCNmcJZ/6d+S/VhyXKTezhtltFeM
GpB/bV3eXgby+FTEGM2+0eFkHCDDCeUnAgeshs8wK7+8JSZeM3D9ce2YrZmp0XJR6BQwLtLp9CG9
LfqskBwLc0yUHZ1xDiInnSQMuOk8sN9gA+J3jAVDmvYSSibWnnZsK8MR6NnozUMNVgsMMFUWmR4k
7vdFTXD9ZTxYanTiJ9Q2kr5st67Y/UNAR1drG/OqCiMTHo8k7SKO5bhcnfkCYxuloSbSE8QEriUJ
e92l7Qxa15vSIYOnai7evd9KUbdTB02Jfyy3HZIgOJBQuRngcq3UnBBBRu0r5yELvra2SUXD9wjB
suDRxhJGu8VgjsaEOr6685LcjboHkZUc+iQZRoVGxaIIqCEiJNsFwHoNo3R6h9gFnrOjSMoEWM6w
jOaiZ0WYZx5WdpDD9d6s5ZRBXYDLz5w0kke7VQU4OcLm7vWJXLZxoHyeu/DvNtpAtt/bVUj6p05Y
yz/YeEpakLzjAOobAd085vi5UQSMDCi4qeWHUhAe4FF2wgN1Opx3eeZ5d9/6OGvVdJIu6Q4pFrer
XJhcTx+VAwoAZu8YsBbjLwZrJ6l16NVDaMcFk/6/byrNKTqkPB3CHKLtNfIMq0XYeExrtoIaxWfX
L/bsOjrJztCuXZiLzmmaXesUkX6U1KI2SjyFcv39GlG9Aj3TMIxIaGTVQnyyDxgA6YoPY1HUb9dh
UldJFMoEpGjx8ld2H/ZACi5evOcfM+F0nhlPl/J5341+okzAYhuslcP5+iofjsl7nv4hQpXhziIF
gyu5Tsfxum4aZbNon7l+yjH7Uo7ckwFjT1+DiwVlezHZASHENasZoGPocTOCW2iaa/i9MQ3J3dAy
jsgE2fbGweLw9d0cD1uZQq/CE7/CITZuBdjnYhg7OVYSgteuLtn9TCXO03xlxk21Eky4hJm87p7A
u84nya6ySi3urQahaUNxV+vFjOJXB6YOUCrOEGvAhQUu16awGoiftJKiKIMaNT2hsSyqhL025OJM
UwbZXxPc2RUVoVKLtSplWfWbgjGQS1OHVYaxr/Il5TOGqQkfiVH74/+i6bL8IH2hjIBDcoHZbR68
X4iCN/8jvkMZb8S9tfltMba13Dm/tHDzQ/C4fussXAPD5DYySBnzTI+3wI/vgNCWaU4CT+Ccwu1b
aGw4MdhfQ6DN0ERgtpFuyg5yCxGkbts/neepECvdrZWhrS/Pbr/jf4d3FvuEvU/bDXgB706oX/q5
pFwaYCe/gJ9F9Np33PivFJhg+ebZ5w7K/KYwg9DRTnq4l/61o5dZiJYpIyrzkyzQ0o2i2NPvV6AS
CH1O7JUncTkuIOMFsniViq2ECfATg65/Yrgee97zV9QsuAgOg3NBtbNLnQ38aGVpot7oQfGvTONC
r3GH9Zue6844BotIErNUR6Li4ZJ0EsDx0yu6Nlm0lkpCXMeqdcQ0zL0ajXh2M9Z3BbMUQdCin+u8
De381TK3KmymUgb6Rz1SlDRlp+7U1FwiSVgomnjAohnPImFcOVeJF0Wz7bubLTvgETYUqK2z2vIm
jl3GYFEnmbaEdtYZ1mYnIe893JAyBee0dxORuxVX1+8/LW4In3QEA4Ek5d+GJtNmePWGTMxI5TpY
tYIRPW5lYmqhnwWCmiHjwse6Yk8XPekEnstayLBMXCpf6eK0L30GMu3MzpVsRwoA4H9Yg2PPGKLO
wNwEIyjdF8XgTdThb4/VPf9DDYY4em++5kn/SC7MaWCNsST8gWJtEP5PxFrkp0EoaF4J+P7DTNgB
LbOkStpUJrbsRLXSsIPd0+H91edSntROTGguClM+dfmIgvkgioVEC6o/EP1GQLH9upxU/cfioOjv
SOp8BB43/G9kszAGTOArHTodXGzLe5THDKGRevpYIY9ECTEW1ec1ePKF2biFlZcI4Sl5kiXPHTtT
Dz9DsI2tPsYk/Y+ywgXxDSFaMGrd0PziRlQ8QTXCxOWqsrUkajZp83oU5X3lD9mx5EJSrGc6gjIu
IlYBrOTQEDmlr62kyq5dQK2pGjbYW92Z7Tl2Dch3Jv1KIQO7YKgIXYtCW2LyWzbyvxsZf/ZR/5Y0
xjk5Bptv5susNPeu3pNxB9xAsJqALwb9ie2D/3mcbh8y9m4oCxtA919Fi4OotPVDqiX5J/D6DAdW
/0Nd3t5w1msqpyEQqn9zkqh2pEofKsVCc1veTOVzGfP/Try5UqMBUeE5yLtkq5fGIsLzUBMyqD9R
sKeJWfzj+XmbEOJnhSlxqfqQZt8PEInjmAkTgrCDo4LH0loytggHulV9G8H37bBRPdcstP4rkDTc
SDHkHKEKM5RaQzhUScRUuJqEs358360PVbO1XCL3F664e0b195iOTthpPmwR9MSo4aNI0cYjur7B
qsyiDWLBJc0tRCJBIMYq1FW0IrMKaFwWhRfycArwPQbRgALEUhh9LE7fXnN+Q3Pi414V4MVCOkMy
K8c1j9Ky4mZb0CvVIOLG+lig+I3hfUD3ubXm9qg8U3BdoKzItrCvj3Cyoyb/3nVxoJyTUpNWmOrL
JXZvP/yqYXZU2yXikSV6gfggbwvOi2F8I0jSRuwaCZwhQ3YlKbVBveFVlZwBC+LEwWbXBsDlmYRC
I5UfMYN0QLm49XjleNZYbyo5ELYV1nVufVVtDpl/ie9RgUnWPqf6cOy1ohfjoRYU3iX0SU9INcBa
33ODL2OGIiKOQbuksVEOBv4hVD5BNhXhFdG5FsZmPxFjLeDMpHkOS51nxWXDW+w/4yAeCIV/jXrl
LINXmKHeqwHT1Xzs3psqcb34f1lXjvDeaKVaJq31fyn7Nakv7x7FWqAdHsfjWnJY1reUDzGoJCun
adAJ0Jg8iVzeYgbp6kGa/atedQF+91BM5RB8mJ6mWGFzgQNBxD4RLoJsn3aniRPCfPPLKmEieZDr
2qXpE0hLeZiX/Mprl/fhjRjpHrsUK4aVxzT3wQ/E+4U2aDbdYEvVu5xMUAR4o+2NHCz1EV7Z+b51
UOUFOYZFtsfrWMugUomqBLAvuSEtj52IMOYoTY1RbQUcyCxNMyTgXI5s7AY1KZEgNUXW0CCczcVq
iXz/7NKNGVkF5ypWP7VHm/xZVKIRbWO7+umlaAZdarSGDRIZPm45xe4LryxSl1segfdYfzcnCz7N
Uo7pWomv/1zqLYhZwr6wBzXYgWp8WKPLvrlL/mGOxpHXlO1g4X1GxAham3Hg9PRJ72HpbIOavsYP
WNQpafhy0inknWUoTbHkcu/uq/6nnB7HN+cbtx98sI4tvoFcSFvx3xUzHdyj+RSFDU2yclxh5b8x
tWVcGNLKPQNxhJEmnqaDoV9Ec5Fm3HoGJCAtUn/m5pBNWKevqM+OufhLLe4V/sZzFO6ePt4gRQZk
8DK11Bx1nBfhJvnjirhl9jKsUGR9rIG2um/drkuSpJdajT/Sq/SlqA/OVsHlrhMS8A6wbS0aSp0p
EavxP758fxz6hrlBK7YNRmhFZ8q5txSCo9U4XUza8DEIisZ0ojCAPp91jl018iq42vKfPkbEThgp
OtpNgKdy6fsm+Rk+nm2BGK6ri50zOYo95CYKbu9GjILHfUFhXqiWSjKabxlF1d9uJjdfTsoTpvFD
kK3nbxMw5PoY8rj82UDyYk2TbqAAd7vDGQjBSWn3+iRfQr8spbVBtzKzJSGGDLxqfXbgVj4XlKBY
VRxXAD1LVNvrB5ZybsnxJIUIoa/8sG+5Nzp75CQSv3j7jY0PPuUNYi7n56HBIWCzMYiA2njXlTVz
MPQiERFpI/8aywz7jLunNtBxf719cO79WewyhgPbjhs5aUfkkE6fSHkqf9QGnrLVtx75Dttxa8FB
uKG0dCl+ZdZ2IFPJEKhSUNMEJKjBHcdc0al6TSIPOIljPj/HQbAI2XfOJwW254p8ksBN3DTgtWZM
k86wnTVESEkZh4PXmXMqvLIfsdLQq27jfDYVL4K/AhpgBiVNO1hdOUoZtAhKRQtiGPV38vr+zOyD
OMvhj8h2QH8sjsEf+yVNMyJuIIclxI+enc8TdXvUMRaFHYDkiI71iI51az9zcLrmPHGYX2DibRkq
j9cbpZM39AcsU8yZFP4Ns8GjDT/yrcfaVElTiMEgUogsjhvFIQAsFhnSNf7715xm2eNBB8hKaFI7
TeMfUXiHHNNyCgM2iy2k1yfAvMuU1d3flFdY7k/A5ZMAtsxWxJhcD+4Ae5QFKP2ErL0XLL5aGbCs
ogNLgMlCyUN+hVEt5O0DOGxRsP2y2vmGgYtotT2jealaVl5OvIoq1k2QG5RqATLGn9wwJisi+/iB
l5VDPBUJzDecGwciBXs/A7zC/nQ/S8A1mhNvq3XIf3EjDKaLQ4rz4gTjKqYIJvCJvH+EbfzNsnYR
rluU2VJdHaPfI7fEGvWRjyuebjZh7mjCRM4zLWUiQnUv07wtNoM35nEKBnFeqWssicLychqnTYXm
kCNc4XdakfEIEONG5eRkQ5qpe4g/lbdHnp39694QkFciJJ5LAegfjZ5lSCZOVmN/+Vhkq928CxN5
pDGpDEqftvAfhZtBxb7V4UNmJBtnbPZKrbRiS7glCVqSOrqnd72AixDE8yx7Ng0+pgQpN3/QsmY5
muC/A1EXWs6v1PMhbUm2wTDQtpBX61bjSXf3Qdd37lrzBxt1I+ayo8rt/aobW7fezWx8Qnf/vOPp
iRQRdZ++KXYfF45fHPM2rPG8R7j5wX/YTEaHtE5oOIL023U31YFJ3sAxEd0NYyT4QqbYKnTdEmpa
64mWeU7t9ToEikPkUZwerzShXdHu3mAiEn+P3fbz6R099RkUGcHmVrZg4B4rf/AuBM5mCFWC/XAw
Et3phhSujiOSoyGJh1X9NQpydhsIqPY7TvT1H+6PRQ5Nbacg7+Hz6bYgJ5j7RHR/+qkXBVkb/A6b
EzUMwGDow4SbYc4cTzr/O3PSwZqcWUG99C77oCITe5UTX55PR6JkySjYHBvRp9FvOJJKHG7m5lWB
+FRYWhg+dQh7eFbI15ZZ/lW+LyF0TWAArYoniL5AflYpbIxsJCgtiPuP6sTdZC/fCaYF/ZTe94nG
ZM/uOJDQvDg1nZrQ8qnPOsnJleajr5PE8WbaU0bqcE5dBVQAYD4DM9CU70EUiVcDVu4QbACAOo0f
S5Bv0EWGBhETM/O/SMh4sZvJE/fn0DUT7ePzd/fJE7iiM1Osj/gu2vK5iG8NWmNV/c2trGNRA580
2AgJV4OOXgog1/zAB0wxtjXBH41QAAGipUB6kP1mRFQt7VDeCi3Elxl4U1DWFjN2fgV11UJZnuez
fH0Cj7w8ziJMosTcP/QPkVgteYiY/d2U2cg97CBFMESCw+hfZhAPE7h+kMxWbNSmg9GVVTXYVMM3
VB2IkJeT00uJnHmmLu7+hGELlpO6ngdJyreAD1sRRBHLbLt8kOV0+xQH6Uk4ebajwK0MfCfNrQ7z
mSwBARTHGuRFIBr4p/qkugL7/y+G1mO5/3Z8O4nerLsUihoh54nraQ7Dx9MnOTHOfVuPyjkW5lEP
NNLmIVlHccq7Wb5HqhdvXJGKv65EIbqcpz3o4BDPnu88otW5XZR6oDoncA762hOxPwkYJTsFhNee
w7f6PqHekAXYu8sV+b1049d7P0opjEICmMQ2A+CXCKHHCG59iOU2PY5J452Zh8Xq6DT0y2ZO+Zqd
di89hyl9RNE1YPiKrZpbQV7GF18QcN+o2dXBKqE12veQCgsTzZkaX5GiFNUFLu9auji/q19sL18P
Zs4ei+8w17TfUS/n6bWmFM0tKbj6CsMyY1XrVk4KramFSElJEQrMgQi6qs+k5awivVGJ9cu5G7Cb
avdciDX99GMS+tI113hwy36tWxsaS/LM3+a3ZsZdhkEzdzeZXdIybXQ97hsde9M92bgf6Ltcq1fZ
owGH2bHS/4gH7Lm+Vwdr4AzlVxPNncL8RRvlWf2V8AXMaCJmIsmduKto3FT8XrdG03dYeOI+FPGP
/fFhq/swZXEgP2yUxxtkrm3tmXcji/Nl5F+uQ4LbHDjA+J/c4By+FDzcBtuZyePNfo72ARfN0O3B
g0U0nGCjihosCUMwmdeZxd9nCOgD3j/I1B24byAwE5rtSZ1/HbTe2QSDOPMHqOGuB0ml+bKKoDTO
/+tbY79DRownlLBhevqE/4c/UI2dCLzRsBNh5Yd2x4TKXlKMD8kXUP9XIfZvFf9yqZczJw9jbRjF
ofdrOzQhJN7PEduEkCqrLdgsMgOV2J0wH1BREetIVhzy5dK6xJfeuPq4zVwYHezDPTXmlS8l5Qp9
M4r/dnK7oGREVxZdudDBavRozTLDmjynHjxKgPsu1Sj6ztx+SZ+vt106KlSzqRV9bm+unZiq8KHw
+3tn4Wm7wk4P5DJArs3jj6bOtLt056Td5L2QQBQ5yFXTQ1sPqTEuDbSbJuTV0mxUfuz5LGDU9uDc
slG6rqx0FQNDBPK4hQnKssdzYnKjIKytlabYICJq7Cpv3HRaI9p1/SarBJvIfRoVbUoT9iv3QeWM
MkuJD84vy5h6miucsHClUcPpVuP1RqloCuj/hgykrAiI9TC9mbl0quhZIvTC8dgMHCidU4naxCum
A474kHOceO1T89N6sT7ZSQr0BdV2OymsFndGhgfXzI/j2k78hZ+wHLfDkiISiBi3za5BSp4vD2j5
YmOj4fcuNVk2KtUYfNF6+rbfSqHCIszNH/ev/flJ0ZnOB5b6ARJ7eCZ/0HXYf9prwQPY4d9eac0k
oldzM+NAyN7HdqHh2zL0Lj229YBhS4y9o2LifNZSmD2WPwF8zJMkEnAX5ApToCoscFbfj/tEtf6x
SwEtVUxjBiNiOD8bmiDdKzKEpTWZxTzcCqG/vUWPHMkBg1ZvFku/ikr6ewTz/gY0/HA5T2na3lXx
hHl6j5JlqPa0+qRU7D1CwTO8eNmGzA7ITvw1hOjI87Gsby1pT51nHev6cked5H+KGi9rE49x3kjc
hv0/ov1qAIhLE2+Z7xH85diDqLuKe2eUxwMhAJxWUcLWv+nUD4tE2t7WHcMzSWTyJClS/wpIJF8q
U/BMwYtzJLyhwV7cRKpx7C/1Tu4nwYOj5r1pf6jMmv/OFFrCcOUbO8Ob3nMfRSSQve2AMPyB7gj8
l1Oc8Y7YDhSqkqZHcUh7cWOI9cbk3BixvF/j3jKOD1b1L2HKmXHwHlr5GeVBv8oylc+8tD+YeXdv
rHjqfUY85M5Bn3RpoZoXy1TRxflf19PLfq/8Rk7vX9n/UtwFM68HlFGmqlMj0HiRNXKwX9plmY/G
LvxTJutMJoMy6wp/p55ySdoQ/7LTD/WhPpDnXsh5qawu/5uENzbEVGW1Ev8iW4k8j5S39J7iuO5X
eWISoSBuoh/iS9TxoEpNo5ed5oZFYFOKRdhOVkVnIrDvM1hZw6OmGVR2a/onj21L4NYWnF2QV3o5
dH4bokRy0Kn4b9G7CGV2c9VjLAHBMON8Rn9hpaPax5hQ9g9M1uqJD2ieaQzFeViDT7gy1ZB2j5EY
lKCh9iTXWdDSIGxek8dgeV7xugR7RsmMA0S71MdFP9T8peRzZRVNDQUkJsJloxsJCGJYS+lAEmOy
vJlufB/6y/wvJ6CJaX5bYCM/xovhSqWlMVwl0gkM3NYzpzgiML8MQMSboLnv5rU7T4sY7KUCRjlQ
BRpZeLlnDn28essmsgkUFk7w1AYgk4JqBvHmLbp7NmHTIpL3wU2iuxx53PQLdX0ZFHup0iAPTk/f
9+xLt8qZP492ghwzihD/juRMIkaQv9Blaeq6LVW2vFGgHQ9cpDkORGoOvZzI5HcXy6jAJjY2Cx+K
hpmJLFg4gCK/9Obtr0CtWcAE2x18lpu6k6gUn8ZjVksNIQq9o+Q6VE9iWEcJhxqUKsH1BJBQ44C1
aaQA+NVYBIjLrftyCpqIQ1looo4X/fGu6BKorqysffDfV4I/0TuSTvmZsQrtR2WqW750ytHHD6Ad
LBOkA8Ns82PHXMK/+7wn+p3ECrohrIsErfmLD/pmfw3UiJsBwrwATVjJ4DitY8GHQUZQ17rVT9zX
WAmuX4PjNkno4cwGXjeF/vqmz5r9TFeGifexq1C7KOsSxqqOhYitNjRhKOiRyszusELvGfPkLDLi
IKn5H7S94686i8/J2tqPzs+jauAXDoQH09Z3rHA/7IZaiaEYN1UjgZpCcXRdKTXmkfmt/UZLXcTE
o/1jidoJpK8t1cVz8zc1CQ3ICeSF8VL0YXpoA4nDvcqcEN3LmCLfCwTq7fcdMciDTX9XbtoZIVxC
DVgBBQAQ7xcB3BJNzgtuTGlzsjfPj6u3YozYX3EsaPe15BAzz8ysyKx3CQC8Ho1tEoxgKRGMB5ya
EM6+siRvh0bk6UQxHAHU5Vurkqm6/tqV7MuJ5YMHqu7GkXNMwxqNrZvuf23/tX0slS9kpJ4hvK/k
SrbRuAPX9RxIU00PjZRtGZ35JpSBz/wNcVvFdvlXI1ihIfdDPwRh5Xmazxes0P1rgIP+4Itw54Hv
vMmj9AJ+63BR4/3hc+RD0V0QwRJCDEBb5F/M3P4SrfzECtDKpvwyxI4z51GNwdCTDB5tIm8PebE5
cv/TOh0hzQqI4m+zLM+Mr9X8Nd+3qcavNBbkZiGnUUhaCH4iAFIUiZkUvwIC//Iwmb/qR21DfJi7
J0V+MpC0a9KL78egm5M4TQrmajloCAmhz5ZGSxFCXudEmLpwfu4jlEMYAtqNR6ZqWnsUp2XYrJUg
feBk+7Onr0Z+7AXWKAJBwT++Ypruz7Yw2lDWqqUQ7CwsWE+zF4bFN2TUxfNpnvewmyqqCMKVB+My
hH/SSFfxQUTMem9h/2Zc2NkAY023Dao6XfrWHILsLQJkweWnVsAIe6NRcRISSvE8pdz5mol/35Y3
eNyENk0bsXYgUz14fhujxqakiq1VtCg32S6CeEpHGpuaOTZp6FuKpdwHMLMT9QiEMnoAqbC6FSXc
OZSCPYRwtuhtJ+9Sqk0FIlw/fF58eeds+bZQsGTlhyz1yE3YInxQKnaNoOGSbHK/MnN1jAjxhD3X
6c09AI3zmEe95WiLkaSLQNt4lATOaZsBiS4H9JvfkIzvxTkvRT4cEbLsOkspk1/yo3pwC5Pb+bUB
XPEaeL4fPjfCejKKImv7krn/+HK7zxEnMLCmepwKlXGlI9EbJc5woozpXVU9prBE6HTb24voYuJc
RSKXuXnFEaWv112iWc2RNsxC6qSeMHYuHnggBZjhUVfbD5GdAIgFIh+P+FaOfQc0t/W+LZbGC8l+
nIERU4qrgmjRjDkrdSB5cizIvLbYlcA9viSRddWS8jE/UZV9JzlJ0LDQy6phbjbMRRZiZvzHIbT4
QWbfF002zKhytPNuCtceRDCh5Ug7F6D7SGwBayA5OScGvKoT3/U2arBn1pG+wdirm6pH5w+wLnTO
UXHbAyj9eM8/khQHZIb0uTvUF/49hfqwe+GeHX1GFmXyWjk7HcICnfZ++rnnpHlX2lv3khYKQ06e
qPmzg63lFJDL94qGjVeMESfTVraaDia9wLl3PzKOvLy/7Xurzw2TwsL0W315HMhbDSsHAf6qbINO
piuPngORKvoLK9QSxN1aZqROWM+dZm32R3Zr+uRWKL7FqaBNfZpIDFEn96UUNbaS0saBwhdQiJOR
cYbWW1LGIv85KGUsYqlHjIlR2EmzibE8EOdv1QlZhlUp/zDTgcITRoq6c94lXUoSARz1JZHRpc1a
aUrUwI4Spesshr3GjrMIBlVTgVNnz25qhYCqAAeTyHgEJakrB4OdquWAsfbFUQr7tmanjhTBpBq4
aNstvXlkqft4ZMmGYcMwiroAEAf1OcnYJbkMzIssSLoD22OidQgG5OQZTM84h5Sg/l8aqhTNlLJh
L+xmJYd7muPJKsktTVvUoOR4mqNGtwxd+ve7uCmtDb5mRX83/zAtQC823DpewzFoFPf4JSbAgnx5
fNro98wHkTkb+/eWgVmfQQjLxclQQE2bUzrKyfJ2hkkKRGspfPULTK/KilTvWW+BxMSU9ofpexUJ
PNBhVZp7dvz6ApZeb89PElsPvKQo7lsqnVOzDqkPsPX1lneIINRRvwBAKCZdpA5Ie1gEWuDem9bh
l36aHdsGepJu3R8potkSm6tmGtovY8c2if7hFSUysIPjsl6oqK54AmLDjp/TJW3sBbs37WmgU/Ta
KA0i85lK2ZSwNiTnrigTTI26MSB+QK0ag/aDbN7EsPDWLthPmOQnhhVJUdrJBkuZAI4hUow7oiaR
5j/E5u7hKk/ap2fVhQ6o6AfW6R0oY6nxReQiwPfEUGxXI8Y+b/4DyOEGbQzzlKE8pdbO+mFWIVp8
SLPQlb/Vw7+hPpChOMQDCedwrGJMtVcS7ilvvTpyziBZzW0iReUM3rSa85jzmjjLOkABkjN41YlZ
buEoxN5bZEwQw9NWnMXzsV1+InjQ+ehm3xuURAE7gBKeifC6DWnMA+WSdCznRvjlAsuya93r+k8h
J2TziXqdXCbxQSqgTHHqLf3Bclu/YULBJGnhAK2xJKpJW3hezJdGJlZp89uUI1i35Hdqcxr5vnPh
0W4wv21nOyqqXlTCAnIt2Zm7TRX+jgn7xbNCD4Wn6xWGSBuDjYGCVDA9iVzxIcUU0zhpwXjxjfWH
SwH1ysJm2YPihZqUXe6miteeKSbDbycX6Jf4AJWm8GUW6VTW4ek7k0YifdPJmP4GeoimOQcTrKtZ
53JIb2Cw2RJHPMw0gxNdIESOwy2N9Qr7FiBuIXe9QXxfC98WK+KewkdpGlSRpoScKmMLZKQ6PP27
wFmkGnu8iFMIsDQyb2BxR0KY8aZoajjV69kVB3lJHZEnhgaDnTbUtkgVDf5RqWIjDtNBRlhdbCRU
8jkZltRv00RbZLHaq9So8nXt9Bg2cP1k4ftFl90HMAprW0GzaJV7/QEkM8A5yRgXLD7mLHDPahBb
2kCqOc2eqNgizQWMpJ352Zt70W7/RbVNyHKJGb48rV0DCUXMscUtvzAO9tr7PBMRHCJTOIJOz5Re
AWkxEivu55tdc3lSJJMRDvAY+rHpzBYD8xgwAb55aEpHSBH9iFrA7al17wFF7UxDgQErIuP0xzQE
oTmWhs4i6oNz4T3IvZr8gWXqOBa8WkFwf7fbCaylUFljaCe6eTnOVO1GaMC4cujfF1RdjznZLvcI
04ZgTh9hjQu1OpsBP4pVF6vdNnKMWbQyl2ifXJm2J0JWLNKVGnc4hKLMpW9AGk9YZzjb0Z1JgMr/
K7/HPILl7G+IHCJpjz9ZweKM4zzQUMp6fjRNKV/jfq78UCKG49QGCLifCvI1PNcabnlmJHRoWhA+
7MUVmqK+dBH2EW1lLkyhFiSdAIhWUZqWZtmZLW80SP5wfichPVASVVlizDv2IfxnhC3PGzFtk81v
JQR0SEnclUFNEHaJzraW9eFs3qWCHtn74iw1AOG2XOwIqob55lUr1UxKvHiurtx8fmGSDt3+t/pF
a9k2qYcUp/PXZzxNvev4FyhibhTd2XNKB+dga1fjU83ZroYCq91ruGB0EIt3y0fxNSpQGuhDkMLH
OPt1/l2zDindfsy6A6n2lD8+rFNma/LqePLXzDT46dOY2LbNrHHFU0LQSpwBoYjAKsKWyYRcqj8v
mDGtUSoVb/VLPMshuXzZ7TM58jt2ARau7GHOo+IW8LTtfGB7aBKjuVDoqrNlqFFEF7NV1naM/xhA
rSg1TrGRAcEcgz2w8asXnmOoV8x3/43li/ylyE70cIWJbBVlGtlAarZelpWM+MSr60pfkT2lQ1Sp
ysDwy8u7Uaun/HdHHHUucgDQLfij2GdwX5LK1lJ5xrIskvXlg3UM28fRvKwWjE0RO83BtzqftUH0
J/2Gn36a632FHpuQFg2ZbwvPyDMjCZoakPmZPB5TwABD3iN88bMIhlACS8xvdbVGO1iu3R6THyym
TGQILiVS1TFo+xi18cTm3dqzxWb1Oyer+bCHY/d7TdCTVj6FnPSwJ9/jVmqk53VxH/RKsxr71Dzy
Lb2QxtCeFq94P9y5CHeU3/3YsHRWc0t/NuRwqKKX0VBEayHY0/7Qwltf9E3JgjlvusN8qFAowusv
mEYeSTkLNigHckysQuWSTRwUDRUWwoNrbYvdhy+t+cGUNn8vGPvC9Tm7omuEPF3AVHD/pCwrScsW
LqbhMqNmndwsHWf+HGFNNb45iWUW60/QsNgQFtxKnpXylGTwdDFt3eTMuh9cFLza6gPxI/tcpY6t
c4s7EYCp/xfMvhhxuiB06snFrYNff0lFVKnRnYxAHuSA/YwEYWD3aXd/NBDx4AUtVNvGR6SWddR8
ienD8b7fdGJM09lsSH8UucpqiObZhWoM3zIebBeD+gqb9irLk4B1PpmdHvdK+vr+x/8rx2Z4zprE
bJQlSaXgmxftJwj52Fhd4MeKEsNzGBGl8v/eYrtoNzPf7Vk/E9TOaAkPZZp9u9tg3pCNjYNtHrZJ
djIEoXUnVbHWllSYie/OMoCKlHT3fG3aufFropi6tt/Cl2QHifqEXJ60piRy0ANE1kO/oeD+CV2d
w5A5tCqf/+KpA+mgMeN6KbvV59M54fAKUKxlXbaGtqZurUh/OQEd47JQw6SRuZUPvO+9+apbCYKV
R9DHdbDLAJNCERH1qpGDy2CQ4r4aLNtrjlkedHav08jZaaMmXp7hQjNH7vn5rfMu4M5b4n6a/2UH
zdrZpP2wB18IZ2AuHEW4KiiuD+T8RYdwh1s10yZQVtlqRXYc9gOMej8/Qi0Z7JB4uKLk1wqkDavt
xKin7JBB50BNv+u6tqUlhnvJjsq4INFP5qZa9NOKL5IHROnyKRRU0IlW4g9Cpk9B+Jo2vYI1gGUX
zrWYnblKofR/l6Nfkhcf/7sxx7Fo2ZxU719QfrPbXyj9OziicODBs9xPPAHGy3o280bwpWxSZwyL
HYkNgQ0wrXEWIv0dzB2DeVS6gPJkZr0hsmMMXL9QK12Bpr9z/rMPsxf6i6VkDztUQI+hwOtQmFEG
N0Zt6lWemlL4G0di8B47H7Zg7CfDWh+Soda/MgRXmXz29sx2+4ykzcZzwDNdK7RgKQ8pu1FO3Zwz
X18O/65RhynrLZUnoxK6MfgcBGnaRm9k9e+rpHR2QIObUrZMS1PBcnI6ge49a3s9mpZEXcrjDUrg
yfmWb0O0mwTeHuuZLUUxsIeOVHILCbBy9qOZHPfu69Ii/tIYxEcOqtFan+yfC4oRym6/wp0g4z6Z
DoG3NFZHFeWVxmDqCr50JV5kX9eBmUtzFe34ISiKyjixQbv/mT7fUchCOHJt1E42Rq53ONkSrOOV
jIgvRij3rGdc3NHCSdXXiIl5nzF9QEUmLeC6a6QMQeS4pABeTqNirbuadLORkGjM+TS7GgSJLJeb
7yTQH0N6Qy8EYR+bX6VMHj6Sj8bS40fUSKfml3gYPh9IrlykweN8f1x3OGZ3tcCVnfD/A04DfHs5
0Yp7fkd7GakB/zxeyrIlVtV5K/yR7ejsWjoy+J3Bd/Fl5qfBZQNU229yGfbmt9dpA1qsmRpBzd/4
LcbTFew7K3ho9CsFRU1h+AHLjB7CywyY6RoZbr/HvMEI5ySE8uTlu26Z2GFgNnSNLwNwF3vQ1o25
IezXvMJ4KbUFI60xRNeEwfk7Qj7mjdAS2wFi2//brFbBh4HsfJMZ2hGSZcaY0ru+BZ7Hdho59JDC
sm5nRnqvVKSJ4MmaALCtr64lbE5fiR/nqPh2UQ/K+zGTvX2Kjz1FNyBYk+m1kheuinlCrutd7p/Z
bznbRUiYNk6A76r2lsJ+eZWiR+9F2ird8hl7QbAUoS0XPT8hNr9G8rgHG86ptrK8wOeVVEyd4Biw
I323o6y2aPp40FjXMnO6Z7pS/WcTl442RyD1G8mxOY3cKvPkfi+TT6qWvvCgAadcFBJnY1RXGnkT
rZObKVXlr7HgCVe/R8LQXQaLreXSeisTqIPo+aNf22253rap08R3M6X9F/H94qj7yRJuNxxHj7S5
X7d8s621pbkhGHmBzl/N0fKx/++Cz+zjsZCmO3997rNxHK+uoHTI3pA7tFln78RjiYw8tEkDG2ET
nCt6cdghDzhRTB6B+f3yOAWCfvsP9xp+pwz0pZclhFDBrb4zfVOv6LYnE5AzZP9x+wV981SbSArP
CPQQ3hL5jcDKWcZYY1ByvdVmczpaTKIhV9QdIgrKHRwAGOKQgNDvZTbSt6beL7RMBOEAJorRDL2H
GtWUM1nw2hXfjzd24Csmqahd1MdQSAnx9MyIE1bi92E5u+u050BZUMg2Qh7AO7LngurcdJrLFDeW
jtjoweaXY8z77/9Jd5NiVtavRwQXgJUdl8zUVcOHP1wARgzcNdHui7oB/hMyAU97JGdp9kf6zGBp
75SclIeYXROle4z7mpUFdjdy2R0/QrCrLhqTqbXA6FBVKqAu3rYtV0fqlsD/4kgGRQia3DtjU7cZ
499aMiuRvWimBJS3qXuetXVH00NTj/8Nv+ChsJbE+aKI79M7unI3bbB6pxnyHedDsi/nrqP6mPMR
+lG+zbUAeZBRyBKRKU5GIC5N8/x76HEbQt7EhsdjrCp8rKvmtvt/SZIn6gPC8mz4d4yq4Ov8ZUAz
npYcHWF4lb+8SgTfU/tPucLaXnaXqkb0D/68lNYs0TQglOxAffZODKaQCC/VL0HAwPUOsi9YRq3U
/Jxo7taITFiPo8/vJ4xk/rHnwUqV440xjdWBhIgWufMB7Yx12IoGkYC1Hh3VMshrT3J04Jtkmp6U
aH9gmd/zEIj1RtnKDABqGQnAdimwikkBMhPdAAFCcDP/G4dybgFPsodGBsE5bowM1S61rY9/uv4l
T02w99u1qDtdFhvrHMnxDYz1Q1eKE7Gi2rtQML1s4+VFRZKjkxOxAccRl+UQkViewYz1m3EL5UlB
omlC66sJKOm8sRGDvqPIVGmbSKDtsx5g5TRkB6lsNYNxqN4cyZ4lkqB8TCWUxs2e264YTQBgq49E
BScQ49yOT/pFBcWV72fc9K/kEkLpBaQ+R5BTv+1Zc1UAggVOsM2aEYasf+Q6u59jIR7wGJ9jz3x9
b8qKHgkYQZq4WJQ76viu/AmT39RjT+lU9puySiJvg0OOuM4aoIksQpBa0x77zzu4cFY/7Ux3gxdf
N//AbPJrDbF5IOC8dFXlbEqbBZWct9rCl7zpE8NcCYxdX/FLJYNubzbEvVbSna7Waf0iet0z5bw+
y3VzDzK9NRKUbzEPTRkKNR2oN20h80g9/DMWasUKBlcWy5aEkJtQjb+jHKWugsu8/Bf4VFW0jthe
sQx49YvZfTvhq+vi4V3odxL1ch8zvttF4A59ZXHmOOoINmyQZO3Kr/JRSbbEYroc3SoNcgqOKvLc
+2x2uytMPtPLqGXSMzbeK1RvdGBp7JEKKytzwjpsVkrDroSIszWBXI1wrdMQU1JypP5No7I/qont
WX5bQMT3yWOl26zd6uHinH3EEqdIMAw4mR9ZztttqXDPEM4Ito1RDeFJkYnYW1MjoDJy0kqfl83a
nrvu751g961VdMzWim9kMo4PdvUBgl0rugT0Z2yga76WFLqhP2U2zQThR+kilAIwNilBiSqSwTzH
QsHEmeBiPjr5yCled3nTKQAOO+5i5cnx5DTQ/kITf12JCDAsQP+EB4A/5Tgr5qPxE17QelfQI44N
TRs4WtRLHfeVfAEieH1kXgCeX57moSkPwSApu7r9cahOlfYpUhvbH7+yUirDjOvzYM+orKWOh/Fu
EamrxN2Qu8yZ5pTu2QqPuvWti9q0AQB80McCF2VYdzj13WneTo7fejusPL815uTjxsvGt5JfIjx+
JC51p/G+YtWUuaWNPb8fOYq4WLIMu0b/2mZMZ1jc/JSWESc5i0kN4k+FHaL9vwNU05F4OkL8dYES
SPj7A7dkgz6Q4KDStxfOOddCl9FhU/RiIYK/UpjyWsnaB3UpvhgIpoPU2A1XPyE8dh2UUlYsLm7G
O/qPlw95BC4HjjBZmS8egjFPJ+Lz6r/jhW0ChMqypwrAPYpo1cTerKWkNE3qpB85n7a6HmlbjxyN
0vHP/KcUX/WO+kQWjffyZSrMPHb4LxspViZQPCG8zRL8QyetKQPSqbgKdpLnQV0f/X2D6Mr8MF5l
fWnB/Nblp8RXO/xTNqHDTs0f2HkRySSOwdJ2X3kef5xoos6GyWaTBhfsnXhHk/ektVJYsqrDDRZ4
zSKUstanPsjwyWGd9sl2OaEi76kpaW0NCgsZgUGak9DyAYf/E54wdVS1ATexHjW2ZYZf1iw5G857
K0haq40/RvDzAJKYYkbKzUF0M1K10LQLFvHopPQ9aohmYdCgp1RyCTDAHJoOylcMsrlcf8wEUlrF
rPa9vw61NQi3TXEMa8RinqNAioSTDG4PkCMYSgjGwkHs4qPzsPEmmeUOAFgAfEEG4miaVXX9yBdu
MCUZpuTXyeNeVCPWtcw8FcPSonhbhHm7rv4WPBkvXUfDxFZLxVudpuEuDPP5jYR3M8FMJa181iQs
iKgFygHibJ+ZI6svtL9rhjEqPewR4RWL2RSgyug4fDit3XYQcXEp4Ou5nr3O3QZ3NtoU9CwB3oHA
bXHaPFlgJNDTUelYV8v/xxC6E1qnaQqyTJcWTbRhJdlYF3akWHcT5zXuXbsz5jEKWBceAVoVOU6x
JGtQiyEg3LXU2U60aa7tG33ozFhauZ25MUrM/e4UTxOtznbQhfxpC1Ke5LzqyxqGTM9D1Pt/oNj5
9NK2Y1XoAhHR91qsDIsumZcBCMNIOoRSDYKI9Pm8kH6jRjTFIYR/+okJK1Y7L7Mxe5XPsd0FrZ3F
+hEsQiS+OhY14+G6MEUMYZXtS+NPkSOVWPJZAf6c4buWHniM1LRmuj5WynyEy6mPIFMgvnwhE2G1
QolHcFboHHAXybzRPYI8lqIBAdQ2nqAxkBzRxwdXxrouZL6bfGMSMZiFKRFCHrw6CR1GEQAi2ooU
vZUf0KrW+4Kdx/TRMX05w/QTCmV6xTB7Mrn1tFHkZWrzGFrojUdvoHSmL9iIVWsWYxzmnnpqqhh9
A/NyLiwDq2yVcQjSgkNIec6DPmvd3a3OaIQMr6UoDY60sQwcStLqgQE30GXsAUWWAh7CDRIPxCJ9
bTcS7jY+0Rsoe4K4K0sZ/hb5KJ5gE50weuXTL7BJYnnIxVA65Vr+tuS4KiV67yppJVYO3z41zckw
i85JsRZ9noxvg3tY4fcqaUCiNkqRd+cdFzBX+jqfoTIJixskYjVL0MizaVA/o7UDwqzZk396rh9q
Q1ABVcBQIklmgZREudjJyrYwMN3PqgodU1dmIBcVuJP2/PvnVHrEWy390KMUv8KXlAmSCMgo1MH6
2heBFJs/fgv+cj/CGDSLpL0goJSSzpQsz1GY5mxDc7pDuV12wF4IJnMd8ZhCvuyah+xpKEOLO9a5
nWZG7TfeU33ZGPtfWKm06G/VbXSUwtPWZDMbBqOx52n4JzvapFrl3F9WWzI93qv60Lx0kdd7oyRF
X4mY7ccu48fBdkNCDVYvmOB4ots0T3B/L+QNHHkKw8Wet2uKA4o/8n2M4orpXZxGT1Rmj/VnDzoh
p3PERbay8MXnhb+mpi0kjmnvRq4ytBqE5FC9q92ypArpZ604gILy/btY0B0vsb4cONgHHzto+JRl
nS7Ec1TA+qNUhoa34kpg29XS2YQ78131VOcAxwWQwWT5zIIBKzkQ388QLwsOv2+mMXxcQT5d+s+O
hgQ24xkXW4JddBOfbziVsiKMjcH9GJRrKa0VETnHrr/2T2yu70lUaSPPFizqeoa0u25k44XI5xgn
4Bhf/ZIL7rqMyPUMRvumwJCCkkkJyWRaZRBFU7wAKKn3m6AavXCo+JYHPQTzDmh6szEg1uQGAhXc
tRmBt+2DiBp0jeDPNu6GBNpnQFcYma1NUXvCRWun9juvRAoO0aXvqQfCxPo1bubt1aWRzbbyD/KT
wRsqXZQHyibNlqk2OUpliVQ0k7U3LKeoKv4Se2X33BKl3/BNT7j4SkEDHthUW0JCmQ5bZkZjb2Jp
nhv0716XV0E8jf4p3cIqKDoLU4b67tA0t1ZBChm29Y9B5dTdj0MRcM/T40r4Ks92Eu/ecKZz3TcK
dHahIzIc4myuc3OoelYORLWa1A30pWTg4hP4IH29dqbVhlebnXAMPxQ4Va+QsGyky77RS0xGl3wJ
7hJ3y9XiBNiRDw3CM9iOPGogF3WB5KBySC+FpCv2tShGkpAJlGhV2uJtZDF2ZS1E3MME4NEGI19B
gFGOiYGB+YCci7c9HUiI5QTdp1diiYXRbIVJoOXQJKd1e/6Hyfut1YMqG4XZqgEwqeaOewVISQXu
HLtECDhZel3bGB9lmQYSsTQtW3f+1diswx2UlHmbtFsKyZHZR/NopNxYjoSk+3oPZmTmJq/wxXU0
C6I3w0VPwstRCO55xyidx+mOGIkMI8/6laqF+s4DHtwxgF3ivmzFthmIgCO7rOmTy3/tGcrOH7w3
JE3YMBRDtVTE/CKCjvRTBCFbdFzsC9Gh5j3y05xl3xoOk09S86frcMuiD/ne/8NafvOCGlDXrTsV
GponpmoVcGf1+v5MM82XFCwaHrNg1yNs9D+7uS2E39RWjVonYdw/VmeJg10AWZxsJUir23NKue0o
Vo4gSH4casq1JmjMGI8TZLn1UP4cTRQsQohvHF2R/3HlxAEYHa+LEAvixUYCeObwJbQE/8iq1Klz
zdCKM8c3J4QlNvi1Ba6rUdMP9u7Z6Yoxo/UQpYvt97aQKctZvlnneGu51ehdUMYtsK+7XZ72BjSM
N7Opo3TgjfZDgaPHd+NjirQakG4fEsq5lmS+84W3d8N8smF8jYmc9ZdD8jNyJLOaKGj/Dwu6kSkd
050yKUZKcwB6uO8h0EflvTA4Onikya/XL0zn67iTtLBHwC9BBSMU1ddKIIyj/NBgtKUj8EyD2NVY
cZZ0g0mR4MObRpFhxXFFZJTiGV/b/0uBm/6ZXhXTpONoS0NTZE2r8xAOenOW1h5LgWY5zx9jutDq
xLDkacZp+yDTy7zQUxbFuQwDcMGHtANr+noptv+JIfyXBPYufAW7h0hq4uB3KnHdxWICYKPkkox4
VFAdLCw81DHCgEEr5eZcMi67hfvbxakyHM9TtVJjV9M79Sdcwu8htHOtvZlT/BA+QtZ2rilEWnu1
lJkdb3Z2wGqbLLgUnTHDvVDTrlWWA0Fv3RLuEdNmoFMOvgEyjcjFDHWTX49KEDVKUZ2Ye/boW+Hj
oMwdNAADLeKSimoKQSnVkGml+Bp2EMvUawiH/rvZ7ioAwZDQcqk5+T63TNTstos0oVwqxW5dZ8w7
XrcX6SDKYXmx/cOpDGFpcI5TuBlhEfZTD4hCZjggQ/aN03a4Ok317b/DxURFjDNzS6VNW1q0yZVd
E42CgRQkk56JpVeMYR6v8HS8WaPSkROcdVhKk5NmxiNvfvZ8hBW04nwhwZ9tO5yZ2pg9dlXALZgc
Hd+aBc2sF/elzuHPjvD9kJVXT3cTvm2e/tk95SroOsE/84egyxv8nuX+pji17ZXOhaE2EKSlNKSR
PjSTBY/67SapgLnRPbJWhCk3BSnvwnrz38D6QmoUFY0qV5Mds+LZUm2/jR8BjF8UlG5X5hnA75nA
k6qhSw7gZd+/m3Loq7WJGh1WvfRdbVU1thOGp1/yMenIfvjrhtH8CaVKE/72I4q3ja8Do0hgXalL
DZZl0Up20xBuQH2lDRDTRuY4ARKlupN6H5n6bb2G8+zjLVgbxP1l8z7nhMAfJPKJRQubEHTj1s5A
7QwmUrpPoRqbU7R0byLhlclqCe4kgmLYJyFpOq+pVdcrBWPhYgieUkUdfuatsQIyiPJOkbhZHfM9
wEME8FdO0V/AzToWC1iPfg9ZmVoTFo3PbwDDq1vO9MwKyq1yTlOsSYfONup3t2hRrfiAZ42MGWot
uIiYYK1kn+sx5x/xUleChMI2fdZwwVthLfIxroLiVLLQygTVfUQ+ASzm73F62B3sz1Jd9bBuI/h/
C7+qaym/4fMYcKFlI/cgxkmHzj4/3biy2U6AJ6CyQIwSc4lVcmJKBIQ5t0dHR7PoLVpLyfg97z3R
OL7T/p45+1wuy0tUynqot/311yQAoAo5VR051UfjtojhMlJ7qOwzoXM1DsTz5dNVnwUF0MG/1Cq9
FDNwg0eUzKObpaiVFwpJX3V/bV5eXOTfEe/wru19roO3eoodL97c12kP4qEn+af0wVnuafe0OADr
qNM9cjUdvQKgWrcJISRWVhFzL0F//k1mHbWpRLU7VHtmTAgQzHBIh9gXhGclCg+ZCOeDuch2X/IS
EABbYGFN3Gm6VwecwepNJEdGXjcF+en8hxLh1IPOGZWRU6owOGHOP81DP08qkf0Kb9bYa4BBOBiG
up2X/Qk8SgboiGRrklTdRKS2GCT2B9x17mAfMql5mhm7tWKwssFMI6HdjiVgzTunxsUkobkeERXa
X6BWxhqGTvDgXiA3U1iV/UhMHf2+CrQ3G0Q7ARe2zkidYPVOKRfqJSxCfpSnR2L5vHsonKWgrfA1
nVvILPnpy8TyrFUjt0v5BDN8NS23xWtCO0AbrnnSQFqU5AIb0a7p1saPou7wVYi7EKsdKw/nn7Ln
Odo/YQ5SWeRdyAxeNvye5/WZy7KoJzHW9IkjexjGcaglMJn9cYbuaAz3MSDt3Crz7fNM0m6YDkgD
ko7dJ1AUUlYI2trsuX+G7Bx/RWYdkMzSjpJUhqgS1ZTEhwqfI8I6kzCd0ZIDfLthdKUKJJl3APX7
kHOTg+L4y54k/I8O7KG+wxHtpvKtsD9MHpHgXcsx5+t/uBqoi/pgCruEDvIsU/v/PTBnToEANzIE
whfRSQvqR6sfBByYDrMaw2rZvuXxRQnOrQ8g9SQ3ANU7oZv5oXncpPF8B1w5xARFcTXL+ZgQ3Tsq
2FUtc9fj03jshGY6ffvDQY/vg61VginvtMcC5ruoMfYun3ugt6XtQaXCN+OR0HwkNbeexc6jdvbd
nXUeDWp3Q50ZzAEfFVGcU2WmUSvDJUBSawonQuEQ1cUUQ4vbHXjg2RsxqGkHH2HZEwFwP9AIRjkb
M7QqI9fd68T77huVYPiX1/Snrfpa9ykp5PNC3H/9iT4gbNNQqirkf5gHe/PDL/Bii2D4LxK5If+a
hN+Y5LnaP/p+Ll/oPueTa/yngfwBjlLAIDCy39qlZyLilGcq4teIYvmT/mkQJC1uRvdFoatO2CJw
K/rk9SzZqu6Pn1sA5/fi9kHi4T0yqS6+VL7K5Rky1czvo/N8YR4dq+HHrJus2FPw8QcnOZEe3JtM
MERdSe2x4rWzE0VTmwNRlDDeHgx0VdbwNM8fu43hTr+RJG1WO3r5+4PDtUdCOLVoWvUDDTNEwOFG
qwGOtGlYkpZwiGTXuq2gnrYJhxzbtAcrrv5UXQfP9GTE1LCPtKfBGhyMFIs4tQr5hfKLQj2iQ1/P
vQR8FXBY9fMsJNoBg2d32NMD+8ZP07EcS5OxsCQyH9de8wspjiJ0+eCClXIdGJ4yPaOQyBoWqyWZ
A3zkdJjiKFnJIV0VBWSpaJ8dJFqDMev+KgWiSPw25Fa0zkz9qUuoGAq7WkSOuuqWoe23Xz777B/W
/M5eOI5HmmdaU73/yUP1wfA8hwvM3KsLswzOOPUrGZbLVQgB+CPM78H0jetYYLo04VYoRIPypkad
nTkaSBRWO5JLy62vDjDTK+OgzZMUsgXqIhr7qKo6NhoIjq3GWKSri2LW0NdubS1DVnAuWkvbln+D
ni+lAPSYL29Fx6amSzKqP5asTykkv4gpJGWTP+VVSdMHZZkyLT5NB6ZZAdu9xcBQoCQFLVNIB7vq
zEEVQfuPYtRLYOfvjBb24tkIxp5BCwW01jm4fbEDKRXyxXit68VUYR8BqfJnTZrrUyicdrVm/Cpw
pu8cosguY/pLS0H5nQMXMZcSf4CSqMeZ692tEkTbfoR93OIb3Xm/Rdd6D9Ocv9VB1br23qabXS5D
qO1kytEL0eFvuH8iotUVqzAR/lFCFOl1oy4PrklP8ZxJ8YrRwahAhB+XH+7zFsobf2sPveHD2aSK
U3yF1oHz/sTgd7pkGBGXbr5ZoQZN4CSV9voE72HUtWrNAusRJxWpiFa7aenL7dr73W3kht4vzApo
sogVSx3yNZ+RdUL/cEIfz3nVeygTkZ7FRU4EB7IJtzHoyD49oZEa90EHRX3WAXPI+G/24RD/s7tg
PtlCA1iZ/kEt3Aj+950G8Eup/AQcdRVI6UxIiNx3YK/8GnarCGiPg+wCSsBwk2/alLhJ16vj4SVy
JiRbl2Z2mI688Oq33LRzK8sjD5EX201Dx+BYFo1iVLmz3XPupxzLqGjlYfADuGTcC+zIpufhGQej
ju1is7XvbECD1reNVN5RFOjOtdyQGtAp5OD3plCmVuG0QIz+bmSLi3U1kI+7oMQCRp+JJ36ZfLJa
CdQRC2eEj4Gx+I8TwtHOrlCxlxaJfeRdSXANN4rftHMgIHd6EoxolJ4Dg0TFPLC0GV5i1VlL/f8U
crkpHWdCxsCsy/ujrAjqLMGI7Aqjk3lQem6BsC2DbQ5GjmbS+X3AsOVU/Jgw74F/trL6B/XXtjBx
7rcOqXOSSv4qSbAUwS0ag9eY3794r0SVuj+Sj9tTC+sNHp9Y+se3EOXTlp+a4K9kwUjMA3I089Gt
yLLjJof/UZ0nlXYmRgfAm8epzvfHu1j8vsKrhhxbs8u5YiavAeA/DygccffjPDNsPpKenraBk5F7
TTHanjERunLjrj8YVAdvht8SB3NmNdbEQkOrXGc1xPmWpNNg3CK1IKjNqXQWHwfq3sH+4XolS+JX
KfwkupDWkEDmhdP0/bfmfeSZj3fsvZkcAG/xmCCuNPI4N4jK8MYnHGffJXIPmX9IqCM+bUbq3Zct
vajxvOsYt6CVPXynVTRKwM6cZK+zlU2dohD+PwHaBOf+xt7iC46mF2+2DCpsZLq9dgX5pXs+Vesq
Ym4lot9rAL+gz+LzvclkiY6T2luFkKjtu7zEx1KOTXvFVXeNZdmQv2ga6linc94nyJWIQHkQ+2Yw
/U7sFcYZ7gUsy0W+s5T0C8coIOH7o1vEBuraQJtqORZ7be7u6C50VSen73FCRR7vMxnSkPhb6Xlq
cjZtyYzPKzDZ6qY4B+85EIyDFNlEYxv16RrhMkyiYcJ5jlPHzgmy49ZxnAYK/sO/bJP0OeRda3Un
jX+Yhr6apz67LMxRy912AiqQ5pPwMRFhj8+BPVNWZf8n+k75nPOFMmceYZOZb0K/VQhcU+yvbAIk
ZXviWz4Sag+Dp3ujZYdnpXQQt0kk1puo6rNp/k59XDhVV4nYjmx/idD2mcdjqgKCdwpW1E203cCX
DCfZJWnkK04FLLQ04vymhuf/s6EucTid7MoCUzOeGZ4W3kKgIRUYpdpCHh/lje+51etuVYzwkkfV
Nt2+rHO8NJD2ZhFkgtjEmsNNElC1anPeDRZXSoVjLUHXDruIbPXxA7YJcgeYYLy0ccvj0AMEts7U
rwShl7+3gETXRmMhrKE8Z/z0h5vuBDcehFb1+WUw5Z/SizVrAoi+0YBga88sCFvy2FqaGpTVqufk
LFtptPENW5XTxiwjKd5nTo2srn50mPL18uQJuiCviEXctOvwIIpk5GzYLKn/b/y6GMvXphJuPQ3F
eIR2xbISUs7H3Nqk89QeViUetk26rbQIkaDDuv7rfkFuXFcyOYPG9hRb4Rjb9eoY5zl//wObTItQ
24CEG71aWe2TGkoR3fchs4XrWQCQy+ZM3A8aqq2UBT8HVz+X7cTfAezYCGwdKws+K3+/WdDZvsyP
glL/2Td1MgbDeyNYl1Tb9O3sPVL75+gHPcBRNOarmNktrRMFrcAMzbIksZR2yx4PjsiNo2mrZL8t
IhD8iS3i8ZFU3ba4JnA7aV5+DmLtzVsZDIKE2vEiomXc52BoR3Uf4TSvDDIAQJ5WW9EB+Omhlize
DPI9HdkyUVlKvQBx9Cfo7h+SA8lNDphoLlBOqpP4VLV6nHArPSXTGgGQFk44RAnS287C/phtTW+g
9YsfdinCenaysQhD9uYuQrfqj+aUFJtDQqHon3/TYk8EKpW5tyXfdxcq6b4+vcumcmaU1DwEZHXE
kwBhdwpGaMdbOY0+s9IPxT720yyNGEDAaEbtAfLB5PnVpNbC6VC4Fo6jTXHaOq+sh/lhYJA6PsY1
EOTvbJQtrya4aGr+Nq2qGhTKRTHUtHe77SVXvutUXCjvRhQ2wNhbh3QA9RDoUyLGDMwjY4Zsp9Ct
WX3x9avvmTkq1PNrJrPlx7UV2fC9B9WIWnhMq4s9Lt2GMZ1Q4kgrTH2zJzvqLeucllNcnM5HjuH9
38fyzzsfb2d1r/rVI5/R+ObA0TOd52b4flHFVJzlD/XNwD0FVhz5ggphHDkiKuDi9Fi6dwbD5BMO
mTY1ui94iYRdDrgstlV0IoQBhTcIq5FuEas0qg029ealR7vSwBk8xH/ned1YFtc4IhrBzvx4HWtF
O+ZWGtUJFLrfMf01uQfkAwhhp25ix9xXsjLhmpPq+KnsqC153j5gdjDJkrlc0AcSX8JGIqEB/YRw
TUCkETRb58/vL2kBfKq/VcMMogIZLToKMRQV/CdAAjohMJlCVvpGzJsODVDnoyyOdRTy+KDZP0jk
virU0/8osCgtwzTA004kjlq+3kowR4YWDr+cOUwXRhGxsvIwS2vk73KqMf1WfeucXaGkSeF94M+c
tBe1PsoYUfxV0OKC1LRXx9Me0mZj/XyphqrpnDq+bxHNN2iuW4zg3wPvhrt7p7RiTqM/MSVMnFH/
qZSBDWAsK451QA8dpnAjC16FnXgas56qpcLuosiSJEPD3bsZwdWRrxqNTcU+JeR7BrdyMptgfB+9
gXqqdz0lAK3bRkcHjDt3tnCsOcGqT7pNeKEEKAbh+UcZMWjyZvAdJ9znLFD4K4bgmCBfC96rTFhS
JGxbo2E55RwH0DukdLuu1IEB5hKOB907xr3EhJHFG2bBA2fFpZKYJw7JkInpLZs06OBv4J/W7jkY
ER2apkvdap1wIIyctdcjf9YRkaIK/WKL0HiFmuInaUyWgRLDI9ruxMa1I8tWWwqRbiNf9QHcHzAF
qMUvujtCfaRYa4IwGpN82nsj71hfDW1ilTk41lGUWGQmWcU0Z/GyOVfJsjx67dF+OLH4xjS48cX0
IedOFA4tGx5JqZhVFxv9GKpS3xeMKfG2PTa6hmrCZTgnWmfuR8ZRS9R2bERAapjMCRXWhFgL5Z7l
se1MqezUMzRqNBLkPzeyJjz1t0HNxNVUY6mqRqE148tsnCowneBKAjgYT21WDRCJUbYnWuAvNgmL
QCzKbE0WcALPg8ntCd5rIyPVzjut54Oiw57pN7UcRDD1rKksNdvYE4IldvUI7fMIgkcc0X6aJj6p
L/e1AT/oWmXRGryI9N0xvx2p3dbTRFnNC/7J1lZXHnS6j9daVx42PO1/j0/lG77kAtJCF+jCF8Bg
d2wVm6qnDb3HkpDAmWW+Mu0NfVvwkcqOKW6+ui98NDhATnlWzcKF7LwQ1xnsZXMhCstYn+uvFVj9
G5FdmtQq4lNJJhX5Wwjjo6EkiJiwi8JmWYcPAadOf0YOibNqENpigLoxVcg8RydSsKE9DVmdDCg0
xubwqk9NTXySGKsQqHfZf20cWektf9jwW7e3Hko8e+iKRtChNRSH4SQERzR1Os9dDobFlOJLxZt7
D6Mjn8KKOd2K4u7xZ9nLJO4O/obppPggMPLcLRa3XWXeuhuGGgv7DuI7NtRuLIm4wJ/pJvAKPJuh
XtydV77WSPMLnixNGMmRJ6r3ywAwTukrFD8FYw8fwbo8D2QAO5EFqW7XAOHk36oBp2RepJgtXp2w
vjehPbVrNAfz0TI8AnizrkGgf4YSu7KhWg4RJL5Jj514zx0eYzZ+kthULMyqesVkHQe0rPo7+sGF
D4evkNQDLMWzkAxxOhsoRkAYXT6CoVj5lEvB9vU2Yrc7eKiy0+zjqW3gLHsLpoM3Wvpky5W3pVsF
Cb4ROuvRXhZduaXtcZDmYxnw7A66asrKv0MtvcZS6GbaO2CSz5b9lkzD2usHwa62vtbN8X+NcdWr
Z5xh5/h9Q3CvzTlv7OURpUjpJPDDjvAH5BC26aSPZ8ueB6FYPjqmViJbDLySXf0Wzd+2uhZpqgGR
p3PBcLESFRqgx1uthUF6JjKf8QTaAyfnHpKZDzCMIlOVsGGs6eZRFNCPMRFE4gcrhp3oO9fe7r3t
VYEmBZRV57FTZrVrzEU1Ao0YOGV31NBDvNOY8iLWreZC5mVUKpguGkUqCsUQwNKoUUlxMDBA2Wj8
cULEzQrNCiLJ3nC+EQ5IKokgA8x45uHRlmATWVQybUrEGqDcCXqAaJ2dWLKiLYaY3BQE90PlmSRL
rsgSFnpCNmmnR4l4rtnxUOdqgfbDRoUvAUvQYzqpIDfWQPQAtvWPxo3Vra//jJFYuid0MmpJJr0q
twE9XZjUQcvBBJF1lO0dJsBuKSHHW/am2icGy97GUjRS0c9uTyEYImSjX6/O7wSWMNaAR3QEgC36
OOmaCtVUmAe8b+Bbg/AAe7/5xc5VWBOO89ZW1aRrjVWfWgesQgBKtXVb9Lcva50MJux98QyXgq+w
u2Vkbctpijk8NohXDWSxftp8sXSLTlxLRiolbD42fzJpnGrBMwm7Hpw/DCZiZ6KqcVs7fC+1+kw8
LEalfGcVTF6J4WWQvaLyvmPS5Y2lnuLQH1naZ4cFtuPo9y57PsONxkiQOlc6YhCHUxE1BfhoN4SL
HCd5hJ7pBJ9fQT6YwQrGOswfrAd+yL5/WyFemGLhG86lUedfdXIGfitJEr67gawsDj0wHOLWr39G
upTsf3+7Qh3WI8XE6IOQHkjRMGKac5BNJl2EaIcdZn/yk3MoAlRR+qC3LVbahLbYccbksruUbHA0
QnUXO0XsK30pLD8MtbZkIVJ8lKytSY7TF5n9fOsICbbycSSkpc2haNt3eH58MWuPlS70LfhKFCU1
6ZeYnpO9hmWnwUo3t92pksSqZTUplkodvtZT87th/xYHHluCjkGJ38BCMa/wF0nN/UlLlORBJG1R
SnONjzgYEmXKFIpjfkLwfWka/rhHfrvdcW1CSQDaaNOkUPXqfohsBZTpyF4rIQaUxvNBLOM+sn8z
lqmqpOS1h8x7IVluGgmCXLH81245HO1JPH4KV5jcQDCAbtSHqtE3Bes/yMyBQ5UIeJ5KB582spzc
vAH58BZ/LtPUyeBs4JzWmBisCdHOvm0oy5DRUPdaRihwnYUTCyxTGDrihLTYN5HNHAzvXsjIvjC7
BSeoJV5QsXvkW9tdj/Ca1w/3NujSyFVke1+HIC2e5zljxqFPS8Ghcx4Npofqzou3xoa9S+xPAumG
5JsSupyfuGv27SMDTv49r7xRxBmyPjNUakdjwQREkazPhFKZoZYnvlz14wqCTP5fesMHbyy8z+fJ
QrQNhZUNDWH4DDf6gm1O6/vCrc1UyKw7njGpbazWJS+GXSKX2FuFKuL+KteQvldEsyKAi5gD4r65
wpT40tUbnq+ARkoo6mcR6IWnlw7RE9+Wfyw2FgVFYor6cuXO2wFT5vQK6FTQcypTdlLra5m0sJJy
4z4440zeLsBGQ/WNKw8mH73i5bxpazon8t04gh6K+yASKW7jW64r2ZacVKDQRKuZKceBO0z6AK66
qXGaRwWqlYs0NaI+cNZdAHhI09wwnQQ+a4zjvmRQBjwGa44g6wHCJxRFyprPM28OLOAm9spfRax7
KpOHWJidb7GvY8zw9prEmz3cqzI9rl+RRnAvywaMQ+3Uz6t9q0D8+UzKi+BBwQu8a99nu0MXwmNY
oT1b6Wdq4txK9D2LadJ4uU+bvhThdWdx7aj095REsWS9/fMOZ88Va22AumtL8BMUfZ/dX04invWx
XC7y3r3PO/SkFgWEqoEbsthxCUszkaM4uYQ5Wt0kQzCnqakZUCeecqVa9bzI4fM4glivYzLoQyTv
ueVKW+oC2/oU1KJmutSjz/92nmIDP/j5eFnUMBGOpeOvVJmoMXI61L6pgHw9YxU13gFAVdq4f3TU
+0EBpVE/iKl60ddVDaL2ywgMeDrd4dbC02NlqjPjWiEKaZRVu4WWyAtzPFykC6EAYVIIFgMzfadQ
ECubr3e2r6HFsSabcEy7t53uGwZWqlKQFl/0LTDCfD+YBGWOx2KtKv3yRJygTtbvJ7W2B4eYcvVg
KDAKUTaLM/5OC4AQ0YvPwrU17xR5wYQM4V0uSUVP3WtSRmhF2QaqMYsXIrrOCLcFZXM0zQ7WLX+K
3cadYPODn+i1cyXvFf2CtRhi6sqrEXg4jb/nfhWMJpBC1eonyRn48+3oBLJaFqZzr7XbFje9nqPK
rS5tnckA+MuiF7NVSd/SP6nt8ai+WxoS7qTbxsrTyedxR5rWvZtTLmo9aXlNkPEqhmwja2PGwybk
quSLt+RtviSo0u5vFpQ1SVo/CdTLWComjQtUqBCJ69TuiWB8CnxBWVckwrchraZ1+pNxenO2CA+f
Y+895L1DQEPsrxfPC/Lci6zpEXzaVwGUtVrYtX4EgnBVB9YcqudM2h/30b6OrjjX1tyDO2d4Vd+8
n5Npiy7zWP27E2iI5xaUzZfZ2+uPWm78lgCb8KQqbBv81b6WcTrXt5b5D5oW1BIwGotF9n6XkYO+
WeDr8YSKVyal2vtCyDWc6DsTyMI3Yy/yJHjyi8SRSi11CA030/WhmnT58G55rUZoQI0W67RN6078
em6zieE+zP1zUfjOX6z1Vb1tSJG591e6ESZZDwQ3X6EF4Id1104hzS6IOhFHkZpdvgvFZEUgyNNc
Pw+B6j400+jDh6Enn8EZK7cFvBf0CIypmSdgQGsiFyrhVbNbB/XKFXJfGkVWrpq4Z6t7M/iz5N2U
948wzZ+H5WSJBI5UBClTUG/1Zv3LZgZM7OUOSvFg/3Va9KlgVeY11UctojXE/FhC4Iw2WQ8Jk+hB
dRx5rVexbxv7NI7dnQ3attYxTSD1yWve0zN4GHWEGeIfWZv0vImWZ3VN4S7U0SuoHBhvGTCGFQbA
mVLU1YzsOp75mE9H6B7EyBN0nlCE4QcRDhm1LlngaRp96hNaWQuaebEjUq+992V9cHODHn87A4Kk
1dQhuVJ52iXCjdiJOHR8CJRv/2cdeHHFkPZcJWiZ8DX7De8eSbdQJpIdXZ8l5AGvO+x6ibaRLgED
QxpjkdyG3YmfOvuY5J82W1O7EEbtg5R8n8mptvBz3jiNJnRJqr5+oFfQAtcOPxmjLR1khSyjwqi8
yuaRBoPC//e5Qow6S8fs6VM7IOU7dHPsPLc9elapgEsYEQSNc77oPe6o1UtEnDyJGAf8VwZTOX51
Z8fsrOmZVnreuOvelQbjysNtnwn/H11SaKdI0rmsjXLq5o99vCGgaANYHsLEvvK2cVi/5u+xQ78k
woT1Y+fhZn+bKSxSpuIP1Yo+h4uEDCYi6CepSQLsIjlF4R6vsa4Yh+hMgCWSGHpo2KrEvt/exPuX
r8/HUPoHf8LbYSICgbjjRwdG8Y77Gu3Bp+w4LuOL4oMPRYkAtzNUwA2KQHqZC6Jr07//sVkNnu+b
IGwKTFKtFd/RTeC6GJIcjDkQcKx14BWpw/TcypIT7aK/3/lxGc9Qpzf9e1IVs3dEk0c9gUuUtMWo
PVq+18WFYITuBvB8xPTv0cvIQMaxBo6i9kI1I/G455QaLZfDtQ2u4+MkEe+gT9mnSGXrF6fs52fy
o1/MSipfwDC5CR/fj0KZK5kNmHnuF3dU1GNIG8vX3RGyhJuAifA4p+bpUs7KkXaJHquVLEYRLSy1
ZM7X7ZHYtoCviZkKyfyU4+62ttaY3jgmn1uYDJcY2fp8TuS25E1L3lfhZ2uCfp+Vz4evMfypJZk0
/SElH+xIJUdRX4bbuMqARv7KSMCf2xd/T4QFdFOAriPjdFOgQ9Hn8smhTB517Q9iiCFi8w7pZGf0
EtmH1kbuKNZNT0b1acjQZBZZ7KMFDfrVVfpxYqtbJ9TkgHHOBE4UQ8vxJgVc5/IMHyR1ALoFaydf
uCJPetvasoIsneqeNEtBCvMULQrmWIWSeTC8BKwB4NERwcSqfGhKYw8SYOm6uW/vSVQH76T3wNbv
BCa+fAcBw8lQYwhfOFBPC3qYwCPKnrtCbu8I6v5Lt+2O5Pqb9+kY2JH/q2z7nRlzxXLY+IzqgX8V
Hm7ZQf407uSijeYbV0cC/9WEPZU0BPAqH3gaajVvgSn1xm0zRmxtHf1fCLFdCRzrwhEPVX9Ncs8C
X01yvgZs2EHn8urW6pVwr6kkvdBKd2RcinJrMb6L2vjTS91pc5XpTwAvJnhEt6aOSRreGi5XNinj
KD7Jeb8kER8nA75fd0n1ugza6VsQEk6vpOmBxa9zoAAS7wc6OlHBZ7C+ClO4zV7CjEg/tP6eCAYh
unNz75wZyM7/cd7QfLFcXL8UAmX11WYF+lRHkR40RjnAGzotlC7iAEd8BK3r/rxomIZc7yiYiQOp
glYwl/gP4VZf5jMIO2Xp8FeiuZ/vB5WpgEEqfZRfxN4pLKvU+DZHHoqL7xFKwsclpxnjPcLSYPM6
EcYzx6yG/I7Dh+NKbmYY2u83SNhv3dyxZ2xQB9NjJSsepd8PQpJXjn1fs4C4dTZBQtzL8Aku07nu
T9A0PrY6ZLDBs3ft4S0uxXuvK02r0mOA6MtDTAzA2hTPfO5EcQwxdmRP9Lhv8tXRBh0Enzk/Pneo
J36HyZCySTragEi8EnBV6RgJ94+NXt8A0ZDFuKHHKKmS87g8N/22K+kjcu0cyAoRXr5JHb6y0zi8
LQKAoheekLoegi7P539/anFxwqYJmr20fWZaQ0bVIQLl1/wbEerrIxezAiJBqmKCDyJS+DayQ4h9
Sd/s0fgAGrJamUeeDzmjFo7RY6U8w4zG6AzC+2/aucEBMDRc/R/8TM1t+BUZq4z49e/FbvcVCYsj
9C+F9mnxPDZvRpi7NBZekY2bA8IUNpQIB8IV2mG2OLHc6UxF+DJQJoC6mPdXyQAuvIGOkCwQJ2Fy
eaU+Qoc0WbeNxtbmqm8MeUbCHet6LdADslVZS93m+aMPCl/eM8qaijJUYOABVoYlWqQidSVKel3k
wdCc26ghTX7HWRmrEUFFuAlK+RINLfCSnbcUqC1GWahoz2bdiark9ODUZ8i/FBZNfhRDs6ie4JGp
h3wvZI8LV1WkIR4qvXrkWQ0xx9UkuWiqUR9U2MnAiIQqVtoPbSIz4TWKPb6z+NjrxWeBZfmB0mlx
tW1v7icocjKmYCuBw9hzrh+kKX+GBo1G/xOXhYxunGt4ua/yVTqtklWnsQI7dGZ0MkiOktRPiRsl
GJ5jXiMjY/oS3YNhhhkKe88tlr2anR/beiKHbnntoMPf5jMwfR2UJlHIPIF1uSD272+lBQ5Kjluu
nOy8CNkvtbQFBK2J9cZaXttwbG+p74lB22LzIOcAANY1okAd+noUPvSBsjKo+cLyYIwLYDqtJPc+
1Ofd4V6N/zImj6/WztNjl0BvJC44E3Qoic2mEFQDWbBadtCGX7eZgRxaQVfzsvSFS4+hLs3U6WiF
sMVWT7AptyWhBQUhpaa3LMVTDqLG5nTZvCkGONdOmf39eSQzxMRGcgEXKe/izbjPvdYwF+wIdIfh
1XhwpqaMLWXTfb+/s4C14KCEzjzwKmUk5C0D0Eh3dWr+w3+EZtl0o8pjBKBeEUrk6/1hFND8JmSP
TwqakD/4rTc5MZlMvLMKFWF39mqcrWOCFCQhECHs1oyOa3aMUoFv7meIm2KsE9JGY4OLWe5viZhl
kHT/VoLfCVelu7UAyyts1sRd/8fragulFUM0fK/tor4aMuBYgWVWaHImwu0dBv3+LnnX4V3FL/Sv
gJUKSRjg6bNvWrwRxP8ha1PTVrcPteZlSV4nQYCdK1ytMxFU+L4VjUqSM1nNS+jrBuA6u86n2JnH
QUirLWv3uzyrRR1XaXm5XQZ52igmBijLnpoZakE6syEeHCFOPlPWjU5Cve1W+0kMJEm7nJ76KCJc
0T/t4T6bUp/o/KuLrfCFV1ZGLLT03KGfTKNfxboxjGezynYZjksWfoKNkuWBiIPlkXTIPs/k9cf0
NqgamO1UeG1vcv+Oqp0qUCDpLNuiRNTqpt2v1d8JVb64cqnBIdGr0pmdXwQZnZW72OvWJdRCvWDb
MW2MK6p2pNc3RxJNrThSX2cJ9J7o2P/rgpiE+IPg1s4Bh7PlLqr3Hbi9m9rZjoClvqVcl35zgJk2
HqhNCZ9JQY7Z3Dz7QzxVbBxpEGvOg5XUtwfBxNXPYx6cokWMYmat5SqqsUfGJOO4j4fN/vot8pNS
FvoX3pYnXTyD1Qb2j3C6KzTSs+pkJEGJnKFwhy105jPFOSKYM1bWmEKJlmRR3OvguQTb6rb1uh9L
AngLMlE9YTRMbiwoRZagMfxqm54tj3d33UB54NiHXs4UcAjtb1FEt1BNqIq8/DcamS9fLdwP5m1S
q99/+xL3wil9cteeIXLDznbxF7HnIGy9nKg22FAnU3pm/IrEWyJAliEowt08s4x9LnnTux3XRufp
Qr+EJ5ZkijsGXH4bOr0w23yqDlkyPI+QZLueBYdAT3j8YzyBExEdkK3pcIjzpCqGW0az1ol/fc+W
Nc+avK5HGUAXyjnQ/Njj6sLor2cpdVfbfWH4FxzfEdWd7W9D9yJmBN0yAHovFjIlsgNfWopBxQHI
gmCr3K7IkMySAsDkGQKHbnCkcm4UhYO99eaOAXVrONTj4B0HrYjDNaKeTB8GOUAxTqjuUExEEi59
EBS6EBxH9o/IBBRAyqYSqVCPam5XCrzOfl+Q59RVIVCtTpeXZN5qjkfiaOOObUdFEBRoa3B07xGi
LE4SAvEVWhrKTShd55HDX8rPUjQdVKePMoDQJq+8XJDD7as+6oViRIo0j+OayvmY9hcQ/+mnkesm
q9qvD/2E9Gaf0/FZI1l6q7IrloF/U3+yIedZ5OupeSx9la64DcwOeO2V8WQboplTFpNv3FPcJZFU
qbOHwD0diGPI9p+mcg8aQSvcJJAQGWFaHoOx5aZECV7th6gGf9Cajoxp8eG4NUVIQAuA88HSHCRm
GQtqXtyo8UPK2YV+M4EgE+8cQmwTY62bufl999BcZm7WpqsukcINPvcE6yjJF3gL3MK2a/s7e934
Qcfwj9fLAZUBslwmdEC9iUaNda5NI2ePbqqRMql9N9ZJogOAUAjHeMDu5XC+lzN0ixuJ5eFHN19x
Lh/X85NcRHB7mejO/3QVNwDM6uQ2UTl86yDGe4EGeox/33c7x5TLvML0qRPFmzQ/zD1C7UfS1xCK
A9S8Zx0ZEiRwh3jM2qWLvfqod/WCHnT++zb10b/fiDEqpHDnUfODxLpttccVdF9Ih1SW/rlduAVC
XnQHl7b8qArW75FvHJJZBzQIVvwiJGfChV0hrsk2zlyeSxpSg7wxRrYflcUjFCj7lzTWZVuHrEMP
ci1QrL5jZ/sUJmwvjPDvl32tkz6iJO1qCE7AhdlwNZzl9fXTNNJP5Yjl/dpe8a3D+4Cxtlh+7ZmD
ntxBvRDr59CXruiCM1DccqDb8ZrU0qutXai9qIaJ6FMlKFiZiymGYsqFI/5Srig+SUJ6naOXdvEL
vQX9wtW6yXpEwWG5bxf176WA4SGaQPIJUClVWdgtiRanRw50V2EwM1u+BXN4hZYWy2+kxaBgS+Sx
XaVUMd4oVM7Se3m5ijrjQFaafwACwxtMz8FcQCLHOyIqB05YECSmfDPs3RTQ2aTFYB8pzdLMimH2
LJiEf89wzgYLMtEGdkl7SMLpj5zGP6g8VyiebdIapJFPyyKnFHRLp328o2+B+FslPuF76WGf/FRd
6AIP07Ds65do9B1yb0TF7DZAfr9J9q54xGl0jteqJpRddEBeFZcxfZji7pASTwxofAsvsj8fQtJE
d39dE3IOk2Zf3gKTr4Bgouv2QPaUCGZ3SfFlVB27sjH+OblYvCSQN9CaakBWp8jUnAQz3hV0WFG6
e3X0e+k4rXsgcJGT5PkxHyFuwgje2rttzr0lI6ty9NEmALm9U8r/Qshi8SjPccRnkUkdMUD/3qbT
fFf1Ma+foxUBr9HpuOD4aiyCjD9CPiJZ0hVCVd0EprfQ9PmPzJEXmSXUjX3zcgrMKK52Iq467URz
Nx7dbPcEdxEdd0d51IB9LfA1hxYtk5EDD1xrXIPP3mAj65tGVP93nON1ED+EVCGF/BVgejq6k0kh
CHheUBLPs1J6BUiU9w0ANCRKMRYkFqZAjkR9njDQcNLhMmKX6EEqIbIaHicBy58BazgDw2plwCFF
QIj4BtYwgx7h0uFC+ti1Zobso2MMLHxVItQVPplf0BF3ZulGVlgTKh8PJJyPlh1QoNFIOkaMWUkL
DxwD3ZHjX66yx2eZg3jA2xVx2J97OaRu5UWoswL3cemmS1pZ12sdGofuWyOhFZAO3sty89AlVSDj
vwt+/xIrzT9l7h1wyLSisFxO4gQgeS3UysCCzv9R1ohq/aOfzR3Ee/xKej1I8jeHe89yr8KPMy3i
snRNp8I5oBFDoGwALEM5kTCUvZSv/qB+Lth7zWlFm85BFlCEdaeJZoWrO98WSQv5GENeBN4dBDhw
E2vKkqzqDu3ouFQONpUGyYYJqF0k03Mm4dHVI1qaIKHO2NK4ZHG+xSVqLo9XbV+XIt6d9SOPgaS6
UdqjIAQ6IqUDmR1Qlvj98qfguLqXf+stQ1W3uIkRse5Bh7Dp3w19pgk8Wzivr5wE7yYGRaqhev/o
GaydsaHh33Rw3mhuGyBvQOeANjPdxLINg7Um9vlrsqfebDVEXCmC5a1l44IZtCLh3qHmxmaV45lT
82bhRt4/xdtlsD7T2bWfrepMfNFMqoFu66f1MKCpEp6ZiN6SBZBqcf7dpf+SlWmKZNP7snTEVw+9
F9AaAC9PmaVk6iVvx+JnGQy32+7MdDAYx/qVnf7gJExgYOBrZeRsMP2XQenTFSOJSS901MRZ+rf8
HBuSvCEPWui/HGXrIAFmwBuz+sFbyDHGGbIpqHHQv8fIbuGZmKYGNYsEcIwEnDpdku8b4Gwx99X/
aZPG1FNwl1hpHDc2VM1nL2yo+wHnWP6jfUYyoUYpVpToTL7rTnMSspNfVBUlOOBsy6UD6jnjSz+b
UCEyjfKGU38bn1HkTHx7pt13Dg67v73kdg8Os2izWZh23kZOujQ05Kc5wkVvj3diDROvKhTOQsgu
eTtBMUBJxwyfA3p2QlzX727USZiS6k6rAwict0S/9AR3LWlCISYuQpi+XDX5cWB7x9fuqBmcjl82
XH9itpzAdJsaSlMOgBZg1ttUouObiDzPM5WlaO9/B6CB6vYx9r9ra0atMQeXl3HYwPnop23/th9k
x7+PSYu/BgzuUrIe2qtEyxLYYBqzg25wYViLqNTrbyPZ1SpfFqZSJRiEVluE8S2ukMLY2QTf5c9W
Ir7DKi+IajucsY0R/t1mETwSy8qiSxXSBSYZQ4k8XH9WBV4HTcSfLhL+8/O6QHjPMMXWxaWV9hD4
bPKBds8lDek9kxl/KgPAVtriA66JIwphY4EV9KrfZnZxIQIQ0EaqRwTWZ58MOvN5IbnJAaZjXno9
jyto2qpdgqpXXkWRP6MDrvLRSmcVKuZ+A72LLkObNo51gHfZOCDXA7u+1Cr0EaipLHJpSC28n/Jx
SYojS5ird2Qi4M0vca3IPNIESKQOUp0sSyCqRyOSO/omGEK/dCi6QAfF80IgN0W6E7RiOvUZOIYS
4BBkXl3m4rnP7cwnTnzZGhsgn3q/WZZQdu56wFXoJZl8zbtRg9x47F0G5tNHzQurQeo0OtLZD+iA
0avSjmPafSHr2de1WqHCqHGECuC4bCKn8O7xnaLgW+kF55j6rmUDkV+FPEUjCKBnpSaiPGjkz8qq
bfkEOO3olwVzfZJfGuDwHp1ltxZ2Ttp3JFJsGyhs1tNxciBBw9EUbet8gnaioONOaAXYt/2I0LgO
PMaK+nYNjNO/PssLTPh6TJzVtCk5kjV+TRPghKIW3LUXum+BB1C3lbNDWmb0564ANMLroOisgMxy
LsGm5ENUtmg9k257FECB/AKB14tuzepKmetXD4aAjcrYfuVRwgVsP8lb8879+/htKl8FJnbWOPou
uOZtEA35uM2hfS4KXGcZWwst6+WS7J/4ueC0kOnxAK2XWaIcXGa2WN4ZFu2qwid4Xd6aEy3vvzAK
n0CUzBvOEk2LJ9JTibO5EAqooD6/TDizAQ3xN//dEl2aMaits/XkCZU/+UkNsBmkt8FEqZXq7S3A
ACIvKw1LFK6y8AdXWYEBbWmzRg6+r2k6VzBIp06PkUScokpBaeijfUR0RVt182RgNh5/R5UNAYeJ
3xqGezVMTC7zwoyfWIb4RUubCyeIAASDIcFmAIYBpi1XgJwtYN0pnYhEso/pvVFQ43Q9TxZq7pxo
nwOg+NjdfW+LgZZX+AGXDE3CrmuXMEvsgG/EPSaP/bEYLxQrKUjhFYgWcMesM7ZNRYzmGMehHdm1
elZ243hD+rfrIWw1PRv6BQ0UO/Wbw0HVxngwgrGCvkdKko5M1bxfFDZ2eGWtt2/XA1/K/RyP6i7l
z1qXDD0pQILLz/2S5liFe236W7szFZHOJjg7FSgsfz8Cf7YQkbowYnKUj/MMB0CqFyqKPLMDXQJW
7ZJA2FBtA6bOXHFqIRQxRHXUyTxj5ZnoY7M0IkHoqOmQVFOegmUfbZGZqNUJ4mEHpMa/DN/4iIov
L4MWd6baBVigl13uM0kbBBwIT9aPUtJrZVGex3j5Gbc1eB4m0XPlrpkAjbCccAmiJRcw58pP6aXU
HIYfMzP/3RI3HZ6YI+VGJDnHUBPwpLWqZhC1Fj374G0jIMKdjfK+VqlavqaclLJIiTImIlDxobhg
yE5caKZgtPDz35R+lQrfqZLshw7kMhdFwJf9i1eVw7tVln+cpKlbpyNpw8OJ6vCDA7teqXQS0wCT
Fg1GuRjC4QLSWbZBA064gZlEkzXfp+8DdOyYIcDtEwNcVoWVTZ+LMzAb/LwMikIte7YMo7wwg+NH
jheIfvESFkdC7IAKk7PlrhDPIWASNLxfRYgM4z288fbE1WOKMBVazmfMY0LhBMcQ1W1v38sUtgLZ
9VTsc7mEvNi6hzfWQvBa4TG1CL6RAvPmDwJQTwaDTFQqU6B8Opk4oEtreTfnJiTd/h7AIPII+Qgn
M/s19uNKt/w3MppHToLnf0tGwA8nGzHRu1im1M5Ixie2tqDIt0RPFT7wNoSHE0vUG1vWvPSUly7Z
vyB81cm2kmTy/h++VumMJL6t92jCRRv8VWVzfvPvwp3f0xl5MLJ+6uJqpzkc4ZQDiszXoNexkjI3
IWcG1NWz0mfsbEq9lw3dx7cQJsQom1Uhnd9VFoYZsqG3kLOjAwEjqAnWfEMiv72ky1KnbHwgA1Td
Tk725HgyTxcx7VP91ZLYhbXfDJgX5c3MB2fE8wOF7UHZFMDrqcqY31RHgNL8nvwWlLnyf6We/vO/
aFhht2+6LxYSVtlukt0hS6GcWTGpWKXhn7ioZnj82ZpoQaudRZF9xhMZCTrZ1bBbgWowlW28mtz3
RNXsTQPm1zVPbiX9z8NZRnsOQPcFPhxkpf+UFkL+cB5T9UP5CCdP/cqMTpJAz1dS+0KMBI8PiCgZ
4CWjRGhKIVlAHvTd4mUJGfyEfkvM5fqHgbEChTeH1HhiAR1R5oNbc+x3PxOvzRAxIeFI2YJ3n449
Bu0yvjBuJCyiNqKyeI7vGrg1cvEsNx4d4NyLwBVYeVlRrnjU6/8uLut6iE3zLBNwDPR4oPLpFjNJ
Nj4d/2sdnmvtEsQvuk6vcFcnbb1a7VXdj3QdjquGmXA7SeaRMQM9Sb0BTycFLgxeWH1tKZXwOg/8
XJUEULxWySF/M51sKKWyb/ltPOCDAYazw4FWCKdOonGaocGCmoXVsEtPVqCmri+r0mspBODFzwW8
J0AgO+yYPEWarKLOqoN5iQX7ekLJAFJzeB2wAwnVjM8bXjPaUAsiiozPQBIPK4ruQ4kMdA0+IpPc
hZwV1oqF83s5Imy2elfjHPXP6zvBu+XGlJoOq2VkgdqPqLnmrqZ8Q4XinlYrcemYewS6pIeBjTRz
qOzjcVcIuDyuSAUjf7vCM/0CPe7dngek99XBOZjzU1uOXFTVtbrRQYsT53u4wtapebYErZiq40Pv
p9rcOrAWUvNJA5H/cbLqGh/3PQvL6a2xiyB1m/r2Uy5vIWm7PccqQjc5nWgrBlCPGMNEkKfxy7BH
yu6v/txkzadvuLrb/agAad+eGSPrgy/7wQhvs0tnxN6W+dWl7ZMGjitgUfky0TKVCBG9WgmGfi2W
DX1w96CZf9xlhQROJ+SdMJ8FbIK7DWESyKHfu+VYhILab52BKhvqY8ItHeJznLkPapzQp+eFoGrX
NuY7gTqv/O1y2KqW4Nu30qyFAyIOc1uJsVe9vLPJu7ceHXpxwJehfzngC69VxZMZ+Yrgo16YQ/2X
EPRsYsa3zHbXX+q8BMBcmPqlm5v3FeibZy9+RO8BWYb3b4DXv4OkQ2mCJcCM2wWJtSUv7CBxFNTC
b0ZqB+F7RBJliDi1IfLDXOlX3rZ7VAOUBVza/F8TkljAHHbLT+srzfP+h+HDjB1Gozw0luf9Myd+
hk3NkMeL4BS3jY/A1Pg6rgnsxcMYj3lgXoCwwXWtu4Te9EiB9RLJS2Hxs9y3eMqliT2dXORQONlj
yenhByQ8ESzpRLNwiasRPF93Ti/hewKxZoZXWinjMBNz6Z43ROTg+gXwLxfNT7FP1QfGIrW7L6L9
AKo9junpZWY50o+RKV6zqa1/vfnhgUT4Go1ltoAh04LjnHfSnODvaXZMgeKcm83NZFVuvuG2tCkH
Z9q/8tUTYXLJQxjKjGZzqifQTIAIsJwDA6fHAPbEOLvBtzamUiPFBUSGqOD2oQAQ95X0WkzztosQ
DdY5SN6BS5/A02Nc9ovWdSskdAFmF0nFk4ebktvWWQDxH7CuOSeE8+09TizdeY20WBeaf0jC4Vec
Eb0oHd0wgjXsKK6Qhn1SPI+VhKDRU8JQs2/Hm5eVigPKUdwqpb8Hd002dr7OSPr+P6m63nV8yU4p
DgIhtER3gSuEP3V+sENSXxwcqjuvc1DmFJLkJVuq9ZhNSg98CmwC+7UnxFsXFHxT4oD0Bqbm+Umb
0DNVb3uUHvyA/8BMzIhfw68jElIvkFM6fUdLXB/bTDd9HK5KXPpBFdApV1+LrMiIorMuVLo9RhDB
bdxJeTn2ig0j9w+wfVxlOMHh9W7OjFYxHSoyibstC5911U+cucCAaG7EZdKTvYx97+9sv5g+xCMu
bzRuxgTVlPNzIaS+ICZcads65YjLVp2vcASNdRClTfI1QLQsgSdu0QxUCKfhWTqMiRF1B4c+6IeV
o+fPXuugMpOErr7Z4hjGDoL7TkdQEZzkvVp8YmY+3UykgJjJUu/yOtwGWFlPfReOy4TC1z2P5PEC
PkA01RFWtKcEXEykALyAc3eAyidHBRrZT1wJUqSP+ZeN7ImUEgD6+0DGdoUhGsnSrSi/6m+3fGWz
iQsm/HBqDRgNOpy0hOM0RV8jEQxobYipJzzgllpcwBugl9ry2/8N5+k2q/GoEW3DzKcqziz5HWYb
jt+zFtm5gMbGH3luoUXdW28GIjAkCkwam0ciRCsz8S7xf/H3ZYVAqu0G5OR2SZmcgZFvmsb567cD
NXTsaL2DoK3gFv/lK8pUzmQo2++AmTYAZucl8VhLJKOukQqJ+uA407siu0xoVEhYuSyAtGLSV/v3
4GR1tatcVNuJ95WoDVivlQQRO2NvIbWLoRFON6+1Idh+sVdFQC7nJmAocDRjiM+16STdKevc823L
mFiGJiT01o3V+a4zAlAWgDcI2vYQDTfLAThYPxP2kiKApFCjd2o7PnrRdBocWu5oXGMCrpmY47fD
AvAshYRcEYtgtRsU9pLEe3MpFm7ssyTuGElafocflpHitzpL8slNxAzvRsNwbvHoo28CqQtoZuBg
CC8UigyzXeUHaQFdwLodfP+quiELeGtptp4J6hOOt0QibAniQ8bf2SuWb1Jzgvqdp1J/+OhPMLEd
4NUf5ozZQhg9XB6SX+4guML7fzc3R7o7jMIVgAsZOQ/K0g/RHqxhCUTb6SoV8dmwct5323E6+jv2
uOvtO7OJ9nZxLFRb/odOUGfsvl+vWvcib3u0cP9r2hdA00oXUkgr+yI61hz4o6fj9Uc81R/Do3yw
5m+UsyCgAwVsMZAzhSW2md7JLDkQBs9Qd3KrBXlOEa3PCW42VSMXwqbFIfPzeYarNIn+TuoOgj1S
PnK8p7sJvR+xr0wcFcEGbrxagbxFnv9bTDqsgUF6vd1Y3wYvRmzr73PHB83fqbS6FoSuotrnyr5N
bH7fCZRf0oNT2zKEiapA4GxliPlmZxwwl/kYWJtIsOecMeSHGJblGEjldLnKp1jiT8oxXXACX6cK
MqoRxtAtHiZqnyHdwrHJCKMbmnYvLSUOnBX4YJcJqgdQzJMWhHANDbI19rOra4jAwQx++cma8N5H
OOrudxqxqhwUkOvK5a6pW8NUDAoWLQi/KGFhNctApsokPLUa+L9TMbZDq3albQHKNqc1a0qtARWo
fjtxVChjdAtKjKCvjeVob2mnwtneYvfVhfjU21dIne9tTWbvSzbkZ4nPRVsRktLDwlklWBxch7zN
87Y6Vwhgr9R38vDEmANPAvebY/SkF9Z17MD2yjys+Nt2zOW+8LKl9XyFAv9M1S6uqHFUuISh6lfT
s2UY/tuAzHMKPwLHzjYcDrY8EuHF361knmixeoNgO5wEkJ4W7QYuhJGMg/1p7oTuKrI1dTtSHA9S
CcYAn02uWWHSAxdouFrZR/hWj8x4OKMx+44vT5Nw9upeoVSHMv+vhelTztGSpMzbKp24neSi5zQc
BHbJKt1LMLXcEFh/AX4zrjD9OteIrevf25AFgbmb5K5wnVB+5LHQBLFwn+eR9+fGg7Gy8L5qRjRQ
Pe/tZpNmk2XrEkS6SWaxsLdY8nSnYJuJIt8NtsR5hY5qCzFOlpwt2usJ6pL4EVHufg1+XdE/KNOT
7itvnzYQVvvVl4vogUasrvZ4bZ7J5Ztn/Oo2MErbRH7rGNXzNZX1EtpzTVxlIgQytqyFF+Qdn4y1
MwoEcYmkNU/tMH8oW+eWy2+mwUREFUM01Hgd6LbxzUEIQVkMU5q4eOJA+dYji4or2t1ln2aXfzv4
4wub1q9mN4ahHTLvJ/trubiFa9q4HUyRgnjXAwe87cuax9vTPOE1TAwWLbf60A9uaqTPg1YKh73h
NAkfXh4aVEsIxpDVmolJNo3AW2eYUYo+WU32Y1n9+0BuvVVOAkvOfDIbgR+xR0vDXnBllblntslM
4ZNSkmYp0x/JH/fjfNuMawT4LPkKNaGHw3jNLQoEbtnNM02cyzqiEHJB0tNyzserY200hQwOx7nK
eDkrV9NH0uCNL3gdTT+8rW6KBjGhsUmpL5H3Bcu+T91RazsIS0E562guquRXzzleNzz1rQk1jUWj
vLQweyD25G64qKZIhvVJ3h2zzxVpaOPlMzBE+s+47oO0R5tacrS8IvHfKWs4buWzUyaRnsPgoKml
tUF4NJnJ6bPOaFib1Lk0pKehTTLGjmzl/OZExgQof7jDtPiVRf34AI6dQ49oMA+6nfdgY8l+0Egf
qBKRaSJhgj8Sdvi3PWZwK4d8A9ce6weX/a17lxwBk7Drl+mFxBXxldLXH7Ao3SH85py2JAn/P24e
QHtGKBB/J9Lzop3wso6CfA1IK27vwOT3Zpyma7//I8SwE1OUjSBZr3E0dx3Q8EGc//jVm96DGJvm
etsXIMWhpy8eivo2mfmYCOY7OdsT/kKIRKi7Bn4AsDTX0iLFmgBO4Bm+q43I3lRvMwzeCGhY5Gu7
zHxZN6GtxtbcomqlgF6dB/omw4pTLW68NpQ+DI9o/v+5f6Hsre+iQK5clEE/ziYCGMy2wQQIkLLv
sZJGDH7wKCa0wnjc4dl/JEZkjon6DsCTXpKtwBOkg3zS2PVCCRH7qn9QAh5NJEJ/9MKSqwroP11y
p9/63xd0AZAFTGIUlA5xJWLaceUmdklwKmbjB2a4Dh1Yz7IFmRP9hltjw8dEfTsSRGtZSiJO/+aZ
xgvA/oGYfb2bO3b8hkZtqtpqXKpNXnC9Mn9yF2capZZ0HUKNZeIjW8RqyFUTc3zkCZv+2NNlV1XN
p9vf4AV0vPaLlxNcQQ8pslF4eXO0w8WNCUljy61iOtnWEwjylOR9ph02tMvPTsc8Aabk6SYYuJzj
S2YC3Yx+kh4ZOsqDbboQZRCokyoRKXiv/ikteFZkx3q6JAd03vX2hM8vgRVS6/DZuohVz0e0/gwM
lJmQRdIp5kF6YLYug6nAEbUax7TtSUZ+eENI6pa+DZHDZgIPF+wdkEQXfJEWmOQ+sU7jSfUXl3MS
kvdcj+LCjTgRWqveGZul3h5E0+aj79/mQzPGoFxAY276htXOJ7HdGs1Gy4GezfeAsSjg+Tus90wO
RELi51jeW60M4lWT6YqGV95mdAQHpGGXMzCY/FvG19MFvJYAcHe8TTu6QmJJ6/kJEJywW7pxUtG0
R71llfkAZNKu2bsEjLjNvxDbly/uJjrpq+Spc6MXXfxida18ZbGKfNlGi7rVotZYA8cQm0sQ1Md0
AGRx/22CmVqr67T0KivQE0Y7SrA6QfME+Y9h2dS3fxmmP1Vpj2hmVyvqHdhHLj6pN0LlyCJGH+Bk
TEGihj8K0dEtUlfRuCbFxooqAVpQWCuFW8I389wGGW4kurlqhceZwyQviY5sTTgTcm8ojrnLIqo5
QduggQLG0/cC2/EcelCsDanoS21qgf4WpDhRsh0z0fbyLKeYMS5+breycZ04p2xRW4rj9Dt+uLTl
YtjW9lKyHgf8JIweh14fXi764QLm/Yd+f5RBLdWfn0DqbbO9W7CcwFiPwLDUijk9cdph5PYrHiQi
Xhf58KgRyGme8gaT1DxC1AEae9Q72s8rZPi5ML2rTqD3nhqfrdxe1ajRRJsFV/zRw5W/OjmesDzt
92ti6Y/islkd5y8Nn1k6/CVUXitL7mtqvzi32i1LWC/+Xws8z0N5d2PGj37e5z/2gRQpiZ2OGUiq
R0PMlvARgk8lS9y5UIyQA3UjNI1URfgDVwUd3mU/X/ZbPcN/hCgu+cSp5zmB/kjF0XuAJJnyIBqL
xaZ5aO7W9Hnbu7PzdD66qT5xFC1NkEfTvey8FcmR3Cx0Sl8pwlWXSQpLoKhHcJwoDlqZwgsKwrda
/nU2I15bRgSMAnI9yo2fx51hs2DkaSPCGVPeVl8NT7H45oT4noWWDS1S9QRStJgSacN3EqNFbVbd
1H/qxXmrx3rsyzGXmi3PS0uGnJgCCya/UvvqtsLMHMGj4jujpGqsjj0scVVpJ01hz2K3J4e6gIVb
aWMcjtDj0GUk5V+u/Mzyd+hXAPeImXkzT9PTHrSO/G/iIPuWsHzdi19N35Xy9l/EyFdOihDdXn6V
tQ+uYKXxVDfn9M7lOJlzQIlNJITBgtxdHM62MjRU56R3Z1k0VRrvqqPvGz8odvnfDE4Cp46PyvkY
2yL3I5nxNuWl+AkZ/A4WglXf/x9r/vLWuKXgaKLyEyqHzofuDoW28RzdmIefbrzD7I1KmYN7P6PB
+KqmvNJwlKQ6Pf1EMJKSxXH+KmScvM7cSjSBy3W/9fe5gygYEmjptuY4Gc7FmqeuPUcD5NX89ayR
MrZiWDN8zpGCQoEOLJc3Fz9G14EvTSyi4aqojzPYDzL3w3ImJN0AxRuD1DoJNymNRqxwrhiOE4RW
9BOT8XaTEaakr+GEfxAZKzKoRhv0V4jpSsPID8c8YzglyaWIVwvFGzXSydhAgWyRTZWfWqpZUUZ5
+52Ra9IoIygA3FWO3A/vuNkMCgWdwnz/HLbgbHYh74fkIPb8Ptab8mu3SvKRhhlt8zqxmyrK3Tg6
wqJJIS3F+T9RH3BP1NkoV3kftYjcYKCRAIbuo/wHAhW9L4sRutfnvpH2EtSYg65OTkEsIwb4fSDU
qmAsNKCMkLJsnN2iz3/0RKJXZr5sZu1p0gIiSJvdRIRXNXw1J4mpn29o9xcdUnB/CwnPdQaYfooV
fnMSuUCSl2QFMsNoN4PxsrwZnFdI1vQ/CUAqr/w+1Cfzd6aLwgGCAYePPDCbgs1tqxv7bJlKUrYx
NBZYHrrzcr440qHHkimGLfAnDgjVwr9ZV+7Aaqun4xgvlH77MJWzCQkWDDF4WyOsETpVBKHreKC4
ycCmOikm07FeiTD0Uv2Y0rW9zkjKEiAo5HUQBQW9o96fALLzCI3P8iDimNZ/PWi2MYl/at2mvsfK
UWRtnXCj/NFCz8yAWq03+uAdJcFWsEeWjkE0zEeT8ZMs43nFFsqmZbDOwcRm3kMsTpGdSk2r+VjG
5xuHXsOGnCXYfw51qw4jmd6w3S+g6/Qv4yOjNvEvNOUSVew35c48E14yn9ZPBNMzotcdJNPYqYp1
VNz0Z9A1LTnf2q6AMROE9WcnhPPF9YC2hqUiC1heaYQSAuBlEDMwif6LbwCQGuIZrJmD9DWHYo0h
ouQtHyZJpGfVDSCyDQklmRRiD7O8CFoK72hgPUeyZLbKJ1p+U4IFFoS1WLTKlMYeagC3aWSQMv7L
dE9SdpIiwOJ8/+MoCaCN2+RQDUqkZGwjYf1hcma1Sdy7QtMipeEOlTrq9ig7DUWsc0OE8fcfV6CD
Ctpg0vIaUM+aU58yDG2sV6R7hMNyKsHyLAGA48LWcTKDKdv18zHbHS1+YKl1ejoBeRFl8WOAEihP
IJSOzwpnVZrsxmx2ij/Ftv/Mi7KiErA0x8+1twj1aXTN+u5hGFdsCvVhN1x7jT/vrdw0VmpxurKS
7qgslx434MRmgNPKr8wJUGaawaFWVUvo6/9sRIndtFfkB1cqkQR4FbojKEQm0CIryKKzS7iQYC+o
7lEiAsWapN+6tT2F4brA4hq+MkHxB1LVvLk2SNsnw5ijF4UtlGt610lngtQebV2EV8ZcDYK96A2L
evQ/hp9MLnc7stVHC6FXZWN2Y60xVcf+7YiMsauOjrshGRVT+iSfSJPckhcRfXK+DQPyPHYFLH+x
OXlnMuCxXebT1E3hDBSMpYGGCIeQxyuzhTBEv6tRrOU208U6+jLT+tySO6r8UH8WpH4+fxxWMJuY
CF5Rx9EONhNH21NAcAHscO5dtCduRRNE4FBG4M86rzPJ/RbTqbVNLYa9wt8X+fp1CJWrurSQ8kTy
8gXnK3bpdwOeOIDqeSsexxXRJ6oyg7QwUJ6Ym5mJ19yvzaIhReQNTZXXymYjB6WGsqn6io7+krtm
OBokJAHP0NxwJduq+sKTrLQk6/6yBQCTadbE64ySIX2fBWI7B0cEtF048fquEPfeLUMuFk1BNERJ
c+oyeqSx9qYQkZfACvgnMulCFfD5LWcXfm1FdF+SvzcA3se3e7XqSELidMb3jI44qZqayqxJ+5Z7
UzUYYokrKLP0V/RB2SpmMUZXTrLwNhZabsFAwIucZwHEhMMHJIqioYvjcZwMJSlAU2lOqr8QWfSb
sx6Igi4qFtMse/W02nsyCUBZyI3XeeqGEn2Lr2d2B/BVEHF/6JbRA/Yy1V53ascKMqTYEY0K1R1V
+sPsNwzO0vXQKb1Xbjt2cP+EG52npnBAezMPB04xNhT/ETnZC1vOMGwPJCYU4cpTvfZcuSgxvWU1
1SBK0SCYZ5iT6CIRCw+IpLQBFOmjojekjRQ8sPQ39wIQ6/J0ABfVemt13al3nQCbFBZEAm3qRshq
P0HubGT8vEqkDT3yvd0AECd2Ew5WgJQcah3X+PcRocB3QpoleVeQINl13AjjMdpUFQ52jlrrZe9s
GR7WacUxMwgZP4Zvu0AQ5ETe8QtqaEXIP4+VLWYb6VEACZ2f2O7GkzXvR8LEo5jbngO3CrUkaL0a
TJXlppwfIXixVkF9y6EDW/3q3erPwnnx2YYbHRzS/4gxce7LDjsaSWB2KIq2C38lAhHBXSXsRN5+
l2uuW+EksIj4sXD2SwP24gsNYyqby2XZhLLUUeiRME9XMOLOMYp0IU7uSy0DsHeXEMG5c0KeaU/U
ErTfs4twThqIrVDzVPTZm93UsUWIN0zWzokhRnjpzrjv/9zPQCOmTby1jY8XRqmRnw2G4J2cFGyg
hvoQVYgqgMnGym3pB+5gDX9x1E2TMYOzQxeJBy8w9CIGB81XCXOIff01yrp3WCABlg36s5LzM+WN
+XUibOPEo4lZBeR5HbYYHkz3aNZjPYY4S06yWpwp5OgbgyPEpUDpS005LYAGOHq3a9j4uVttrzCg
x+Q+snNovS+VXmO9NAWAvblanMA5kx+ZzuHjBMdzmDqVNLeptAsWs17uEDAhVk2PKWJlmW+sliOe
zngxkxBiq5YSCrHmY+8Y+Iid/hWT9/yRVLLe6GaeHzds2jEhqFiTyEyt2CEH4aPtn+uxm0x8lE9R
oDtfXcu7z9XtJdSCu2g624Bl1GNEu7CbtkODNePHTQUsc+lq8ITLgRxNHY6ee5/iy/5wksQJPKJt
knlg3w5bXCfyyXVZPd+Kw9V0mFvnXcGXvrHYTVQND8roXu50fkdo5CT9fvhoLCLIStYnqSoc7/lO
8521W2qWYHmowPHQdELcn3AWKuDfhns3Jqjhd+hZAH4Ukv+pAQvvMUmJO2wetsmMpKDXB/6jq2wp
IDOpkOeJqqhhDXecQQaaqmejJys/8+3lQZ3LxzoyK1agKy2XCtfwTQ1cYQgsGUpjHuZZaHs+Sv4U
Ip83zlk2x6GydHOTBIcfkVarXFVM+LEb8l2MrgYVSiJTUUjboi97t7xQtETZCAAZy22dgwOp9JGH
0SQR2D6fBCqvUZBCoAF2MvGkac6PGePcBE4FXPcYeKxctKQ2P+HSYeg0d6U2vaTZiFSuBTzWpy6e
2TLDzgdaIYqIdIlJdHLfZSIoZl+C60sY1dCzAwQt80zfg5DXp8fdheMm9nrDhDYBaglFgLIiNY+Z
eF4XR19sfk+ZgOf+aNq59r+r/q9AIYajDQw2NeluS6iRjUzXHnikW+XgyM9purkJdIEKamPrWxup
WcPC6YoMZnJNX81a2uTMVI/p3xpYKBMsPT2670B/y6Vo0jQM2khfU2+EYgE2+eaZVTCublprgWsx
r+bI7o+O0Li0iLY2HNWtG7ebjH+iBNop3q6PWHQcrQrmn+1YaEXyVmbALrr7iyiXaE5w42Hc/C1F
fr1Yhhm529XZNVfwbHewBw/1+mBQm6TeHEKME/+8Bx+tSrO7WpZjpW9lzxENjhNDrUaOe3IKkTjX
5hgV57xcPidrI00/mH6lx1FcxV3wvLiOGwEOM3DMF5j02kTXYOhWd3qPpF6DI2vHi70C8LJJPX+q
XmXjQ0P0XCxGIhi8j8BCt7zYlxnvd6ztZkYvHgr42rlvFZrN9mKydsRVqMVWt2meNHsWnDhROWtK
/ED37ENjSVGjPgdgG6JxHdEp+swCdneBwHpIdSNHzXuXB15zyjyX2CVD+smUW0GIig+qb+PunZrb
108Y2fieGJjMZlHfaxlVLHE2l2rNLLBOInjpVavN/KZClkL9e2mq+2zWhwfm7hTJzwvVHhCIqeQR
C2WjmadvNsmCaDN9kRmFV8IL5JfhtX78NwoH+2t33d0seTL15FrgH2xt/VZ5IuET+n8mq4x29TF3
BXOsDBNWPfRLwykttX5Avmz9DhmafkNXXUx5a6ihtsOO+XzoJ6KIXZnvvwanQKU6+3x0IqeXeUNl
mjCLGcFkUoTcoGfN4iEmMP7ssLWel7r6ri+fwkBDwDXQ9ozwjIB08IrXPM9jTswjBTN7jmY2Gycj
YqhESvsyfoFdX45uCnsZPy9bH8KDqlu2uZYdbVAlNETGcp9jrWr5YhqlZ+FiELn3IchYnYzGSYpR
rSO44CIpPqNzYWg4ODfygw4+WURV+gLfgg8wcPEOWwU3hoa3o5gnSkSfrWocMyD4FRApVC/DyACY
d3jbMTNst35U3gJRX6rk8s/VUsS+QI79MOnqg34eTIOE1dryA5nDxioprO5NmnjyosbWStpXatfo
OAflSy6NrofD8cEBDPHk1egqWyZrJ5/Q1mNTC4Ri/54YkKNuifRX0ponudxhqO/VAMDuImPRyjBy
jHcA3S4L+NBBh0nK+XUxAju1A/AITiRuntzlZUMP8aWotqRSZxCTFsDZwOUzu6klvxkw3ku/bt6s
+IOqhw3/bgFVHj/+FGbcMNkc7Rk6XMJDwp2YetirP+5lSCkZpwBj4rvsuBcdOliP0VB8b2tDiwad
miGTa/XZHkQjYf4nDesilYygBzwekjABllx/U4Dj0TwZlYLCZ+2yYfQs2AFoTuGNmPPuKBdCaW0P
YQF1dLcUg6N2csBxwJsqOzm6u/TVzkC05MWRiFI6TJdbOJ4638o1UV7xUVuzRBOt5R3ijMCCMYcN
t5+KUMlkPukom026nvDqx5ILez3FgjlzcmZWzrCAlPetPi0jpTMMB/nSD+RmZyZ0pjEu1Tf3gnHq
NbIrfChdO2pMEnwxLp3UXChBzAhHWaUPdWXanyPbRB80GXo8CGC8hti2O9QqEwfDyYYIGp9UwrCe
MZdk3Iy5qhSMtGCXKPwLxNLfj1zW5NUn83hldIybEP3ZlxBzo25kFi0IPeBKvyezZmYAVWW3MT/K
bn9pxUL1hcD3aPCcmpK9+jUfkUQEq7v6B69cBbjvgdjsdncw5paM5YCLPT/L3sJOSFNZW98pYrXL
AUIhDyB/X42OCCOMj0/mBTwon7M/ELBfNMz0ru2E8rVG0u+5HAI0Q3+PJ+k9ZOZb34v/hkPt22nA
jcNXA6WvrFXTBYdoVGRruTxBBiBWg40bl4SVsgusBClex/7NjcrG5g9MR8GV2pR2UOqCz8IGenOO
pD/4iZv+jQkdpDxMrZgRdhrrhJISrcvqITWUEKZTYQTO69oQlwdP6TctqWHAnFcjVHmI3BKyvAMZ
NCPTuEL7WiBbJoz+onle6ch7XSRMamRVZqvvPE4JYO3rQyHFoKNMXXFDsJeEN2zfeRZcBKyA608E
rX9oh7KwvvH0QKei9e4hthx80UVohPFCNn2fGUaPsMk0ymdcsxT3N09G+TrU6yPcot/F/77i73A8
6RKWG27fursfJ7+i7TpGj9rwe2b0pxqeIC+VJBnpOPV54zbgOD4kbTJNE4mXX5a/fG+7jYO03rjz
r+L1M1BsimkiDCDT/d54MGTIzaqJdbWhYztiZbYNzzewIrsy6CqcC9xtwRaDRQdVIY7ZHA9Km2y+
kqHQbLyh+09r7QWqm88NmHvKwTtqkzGMyRbO4nJx9W1Bu1B6sNBklZhNIMjBxM976JlmmH8m8oRm
X1zKsIDbS+6lYeypISWuOw7Z6X8jlKxbIIB8MVVO+g0XbI79oc5lSjQ3LKwYPquoEMW3dPKgXJ7k
dhHdJafsHa0Sz13H6OncKGaN9EDxYxvwU62gjkdSwmkgt46wx4o2Qi7vy6X/NRHI3pWbqvzfAdPz
PXZcat092mRBiIQZTRhJ2EWwJQMJZSVrOoyUowwA4/v2pQoRr7vkdXSAJC/ZelxaDxIJ8D0iNCVc
vLMVFGI65VnAEBS1BxGyczyyLiUlfmwTAXYTObdkgc0qbzoJAGQQZbS7IeuFsTiKztuQnAiWbuba
4OGNd3DDa/utqU+/4h0bOvXr4tDnegFJuOgPNYvwzhj1ar4NFmpkDl5gwp6Tz1ALxA4eUVoDVe0f
KPFcdX0oPrWF1g2zd1VlJ2i5b/O31DUBlHB4txQ5vB9GzerpERExzL1Ie5Nm1s9NzarD70h1IC7N
x9lwfNnhX8+LQIx/WXH0IqGa81s12Mia2mJjUUoYl9kloHoqGPH8Rvj+hLb/D6fLkNF3o9F5XOWX
oI5gWhYOkYmjUsKSgZydohoB0aT1LP/ygNdKa4bjKexJjCAwIqBSg+46uBNMYRb8M6HJEMHI58fg
dV92uMzYsiHkleT1Ra4EMn6XI89gSoXp1rRhqKqq6bvdOU0MxVCSxUzdB8MKh1Xx0iaG4aa1Kp9a
ZiCnIKc2gbPF0eh9r7WJACNc7N8ZAXNJaOoFyfee4Y8Zk82+MEy/SrtDs7l1td5EDREEr0CJhPIX
fYOJ62GlnHmwr32uTxlqIMKA07KkgAsLfHAnvFqCPk0o/cgdZfMHjHuUI0woDGtHgz/O+4n+QPqR
HX0xv+NyfFERUBTSafAw/xrHAn53tfWjWqdWr8bZO/7dfbrHn2fKtcdhVAnX0xCKEgjaIDoWoOtV
j9+3DEmWSypZViRt8wVUk8i+Almh8oz4UYmigDhKAMrchGp8ttKsgKIYiShPVQf7/Usld6gQm0sK
o/nA550+cKvBBP4L9VMp8lPC/U9QyEyjuVBmyhaJBNkrTvmOgu1XDgmID8s16KClNjVdWLNdhu4X
J87eC71BBnXEsaaTrBbIE9KG7jjDbIIlxa9hHmNI5bd4QkWeZlNcgnedJZioFlnYrYBSGdoZj2iz
p0Tc4wf6eqs8MuyHytb4BMOlDa3NHqlNeSlPiubaiQUABDGNp1syxTyZKdGNqd8rR/QUYnLPioDH
IE5KrRoaLbigDhDn4geBf9vwF3XIavlT4Vgzcy1YHD+J6u18tH1V4yIDcYcWPa4MiQTYu9unzqMl
PjXge+Wze0lVUqrhnouC1dWJCWsvOEKU4Of/gDh0o5feIZhaiLDurfHxllcX5MhcgB+/lL53EHpQ
lqRN3Q6e4Ihx/xTdfGmsbjp41MPZMVrca1ja3EtX/PrQXECplYE5fSgYA1VU/GJ+/LxM6syb2kJy
sMQp9/Epew+hXcbqPFIcb+VmHOYjVfr6A1fXAF6P+5+FAakLNM7nLW0MVgmFNk7paaE+C1CTZH7b
Ywfzj0ozQwcZMQLZXQ1IMMBgoQ4ffu+GhCM3/NgBvoV5615NRxOda+Crg47aw+4q8GEEOPa/nvY6
+bO5EgcPT41QeDsmIxlZt09NdzyqpdJuCsBXypUDaSsFBjKVYposWRjSZpcX+ykyEyf1C2vC7tvq
I4a6QaX7MGzUqybNalHoeZERUQtM5ndzR8E80PNy8S66XMYsIgRO5BRf1KscxsdfGR/iFf09MxWo
fr7uon+qiIzwbUa1Hbep4NYDI6Qg2rxDa0LFEtbNZ76P0qfuI2BbQX/21mR+4rXhRLJknEkZLy2j
8bhEXAUAskLGHht9F+JPItVcYKAHm2OGbw1h0VeHwSc1Vt/hEFUEQOBdrXqlx8DiocHuLJkXpyqL
HuhRzKZsQ+wYvZnpj3UbiK92L1GHsavq1OiczPI5u3W3oQA1UwdGAu57Rq7qNN8bxvLtRSq4/Y8N
ObruoBUrj5dBjT6muMVX5jK2o2Q07TwdnHkX9pr1sKieU6B5gLjmw62iYDMfm055DBv1Ma1uz21k
LEhDUMVX2QdVhTjHdPwDbxsCpmKYFBOBukkWaahvpComWjO4LY57JqbUHkY3of/vOYEe4wdkrJnb
1MGRRMSWIHV6uQFSkRkwPSyFLHwfXmNMOar+15G3EUjdTi5CpGa0/xz5sskUFFcpQE+bvpT40zk6
vrujTb/QEfV2rYVNrXTG342Zy3WcL1129IZ9gIKlv1NLWfVPEyeglX3Wtfq7i/JLsQexczXDCI50
nKyLa5VqjfLQgtz8kXzO16zrVgoWstWQWTrKafv51tS1OcUQ8hsCdo/HQm8eTw8jwOoaF7lyCKla
BJv0rtrVj5xWXSbLwXnMfNPFhRsKg8egOYASsWXFb+UWWauGAbYjJrC/JZLVIw1FWcbB0qWl/UtZ
A8aMwDv+VGFi8wTV5AcrIl9Bh75DoyinxR3yeNqPaE92K3PVc03Pcvp/ZGTKTeMFDuxAJAw47m3Q
epz+Mja7u9dmEuXqZcZJl87X93P0DNvjfQS9goL59wWqpKPDqNL01RrtBeJw9NPEyvhTTSmNilCE
laRdCF1lBGLJTcM/cXlPbYdCtvvzq+mKHbL2gRuCRfk0qLIHZl+dRglV3OSqZsEch7NiE0lrQJ4I
SNhqIFCobEc+WVkJDpbm8XZdIWTOH5adqToiy7/hdOcAeBvTeveY8Gb5dtuKMu0oUDF7JYgzDhIu
kNkpXS+hX5H76d29R8D/kAxbruH60LO8BmMNw7nVjMxZ0wugtVUKoF7PiasA8yK+or6kJN0Aajxn
RjGu8AxNWGpWsM4WFhU9jGTtQLdj635Xe/wN+4nInSQI4aYL0BXqoupvHYyp4sixn3FsYEaXIrkS
ohATY3ZJKmkk1YusHRChV3W2nr0GEV78hYjDVbUm/+rJcSog5cfvT41fU5RsTxrTb8OtEP5+3LZe
QKjo4JGqTLt9iDYNJCEZkIDOCKNhOYb2sMAGDAvFsHQtV9Pi3ou0d+WysgQXhnxRUZ+JTA2G4Sns
xMnJQHqBHk6LyXp9L+JXGSF4OYQYvhuQMLZ/ZXWSzGVe5YbHc/vNNFKKLvw0r2g7JX8trMGSFzSY
8SwjXuS51T1ETZlyFrQcfxnygANE9LxTJic6kA/dIX8EjAQugg+DVZVXvz2jxIYAHGQzjcEDxLiH
dindlZAa+uuVeQ8sKoopYV+F4oo/AqoNcoptNLABtfNW27hST1wowPiGjQTcbWNZehnVLtFQHUpM
AujCM6n6R3GzpGqlbB4ynY11pcj2FOk/3UWPtgy2XBLuRekyW2C4nZBB/Hn2a+WzCcH6IpUbYO5M
QoNAOQi7QWrOj+x1Spk97a7rnPZphCkmWpkAuaCwCMp5ebgjVcqEtonLmfAnlMVNmSr7xlEUbJYb
9gmCGEJ3nnnm5/U7zsMewWVed4GSopJOhAcxZYCsoJfL4tb8xu0Zz8NwKjwDl9TlR5DAq8He7C0+
s5pD2cWOfO/1PeYtVTQfNNkveh8KwkptNV0FtmbuRPKf3D2N/nd8O6QbG9YqP/Qo/7WWVzX4muV+
2dM2Ts5yK6LT9tTjsWrHYlMtNtbzJ77lyoYRHzu9wdaIl0nVCx0NQ1dmm2AO7Tz2ZrPRkMCrN3rt
iTLXvWgxWt4TqF9+4nFberkhnvTNOWm07VkVNBLgAXDp0GKqZdpsMZyxAvX24j5aryyuwhJdGvWb
E3Iy6q2978M3XJM+SE7qPA5w1RxToJ5VyjCxmoWDCuhTjseZBT4RMFQFmNNVFl/q0AD9aV0SIwgR
5z/tBKNZOUUfjxDWvNnU8Zr3pVR77sZ6saJCx61gBH9nL+pmqMF5iUF7lRXi3W/pCbsotL9akFjY
YHYVXd1quxOp0yq7NGZYl4bk2P9m+U1NAOX9TyAHTkyqygEPnx7SCbeE9fK+akhCrdN7oKQ+Ul3k
RGRYmW4QBIvBYM/xjlMPIPK31vfO+RLo3DRDLWPaqWxU1HzgQvU1PEjvIGuxL952mZMmX9wiSirY
IcktHkm9ZL1FhcDVsOk2v3ckY3E7f3KwR8c+LpSyNeqeQ3laCW8ZvJWXy8igpR1Ve4lh2Yx7F690
FQHRiClltso4sgx0kEuzS3X/aTkio0GKI264I/1/cCvfr65Qh7TthFjwFFf6m5VCWW8t6rDJ96SH
xlrb9BqL1EXDRVt0PbbT7QOLCBi4WoGW1yMfomh59gaxhchgu5kg/HxNARS6yU0uFVSziCdJeNAs
LNZVVmhtd/3HOJ7l6jG3+whrDtwXdQ3+jB1JjdUuMUlvhTxqa5K+jEkeQXn7cN6NTsbsDhoaMNSy
SSToFWzhCDOKzNVQBzVAyNNglkz1jioa7Tcfr/s9Odj7jI/srQ8sDKghwpzlF0Rf9O6jkwbmKUMi
nkjxCRYoqAjVBRo8VMj3nNw+TZuZ5eKLZZsbxfUroEhmwsc+s5ZjyyFbcsBwn9Kxc+++tJSD9zqc
9bLEslQEweVAKehxMogSHf1T2WpQQaRtL71wvu4qt8aXhuX1MLt819J1daugjRXh9xLExDFkZAqO
Bp2VVhx2mXQgkHQD6KT77da6Mz1+U9Y07/Ram5jcdPlbERB6wkBeF07Z3cCyTbws8iZ1OhWrN3cW
LHUaFDHzhBdHTMtMZFPN8iYliLk6iCd+NfNXsoHqPHWSZzh0YIc4PPnOoLW9+ZtqmuCDlLxUwcov
YBBQp5uFefLb+kn+fq1apO8mqu6Tu0KnopRoTwgLMv47UR95U6Flek+1x4cV4wz1eC/+T0soalB7
thtryl8OnVXLDKjeDiRZPtl6/V9IimFvYUfoMD045SqYEF/J1RXBCzZv/pVez3gEPfnWiZYeCK64
r/xZIQoNovUZU/SzZ1g3BtXRBDXb12yyGqWFU1b3uK0MryhrvtO+yUdGSyaAALpxotmatSeo9g9o
/RF6WdMmfNnjFT7ZNw9yslWoicNjj5yMH/846QoWojikxqKzN9QaXt0bdWEWAfgNk8us/oCmySFH
kgxp7yIuPlXjumBwuM0ZSjb1iCKTx0z0wXjm3rUrUo/XoZDFzuNQkfqmx9PCx59dacdHo0uaZ8WR
0GeLVPoPcrYEVY7GCgR/sf3rsZc2cbrGA2//K7gQC6SYy4Ng11I9NThUmMLaVYfLwPVkY8ogCH4j
zwIQMzt3hfpwMKKxZaZ575nv+Kt7fto+iivMrqEnW0PUO+WCtZpeiaCOXSatrP70w02sDvomFkvY
rN6ioWXYy1r0mFNv4pFF0Gx/zBOJ2f6dLKLU6YBQfV3GG//fFclFgrRRYuPaC9Kkp9v+/5OZD3Y4
tcc9J0R1Ec42fmQQ7rmjmgG2oR++LR+RpYhQSEH7HwdIHoDJ85+8f9lxn4DETxgxg9UU5sbHSSQm
ElqAKUYBCtPlOb6mg9T3k0/GyoKX/Lh9oa9rIiw6nTLFIhGCm5h9tG/KNpgOcycKDYGHTbrypjOn
vLupv7V1uEEBxg090fCWrGavx/CW6xu42/ig4v2f/8HYsQndIHW0ySgQPzY/HgW/JwUVbwHnr5CZ
8kXXwD83P2pcThHmH+6ebyivFhLl6uOsstBUgJLCsZ2H/6+g2jnwEyP8SspsAG+M6dfry654/LOP
uCdCmW8pgg7AqU3tFQrqiM/zrKvfDJBq3KVoI3+SM5yvlAwDBR8yo7GzibT7NmsMnw8UPymXWi0j
924E3gLV8rY/3oKdcUXuQhGiqgL+/Wi5hXnec3RrE1UkT4MddC/oA4K6ACSlNVM7U8p+u8YIcJme
VChqblE3QHpyrDaJ2abmfPXyO7PmkzipWhxdomE6s8QR4FYPzPnF7SnuBR7R0a2Cu9Gu2CcFSgwO
Pp7J5RlZiy7uqrBVsvKRBBknb/UsGbweZlv4jFzjihC0zHXLfEVHKtq2JWIF7w9Das3KBleYi5SH
X6jcbgtMhLT+R9f+jOOdp8u7JaSRF/8a8EcGidgvjY4taD07XVE9W4TVXh++nymTINesT3IlL6mM
tVw30K40gIz28AHx0MW1DEJcClfTBcaDyJQInmk7mkCXOneJcQFRuTnYSyK8C2IrAZ24mAK7GY7H
tHVtkrRqT6vA4unaxiNh0a1QwDm7xhaJuvasfF/UXU9sEtk0F2BV6Ck1/W8ZjrDYbq4FlvbPrm49
A1vyOtVF/wZHbXd3gEOeEa7XB3ZJY4P1iILhZiy7cu22yIkPl760X8B/IQ+sQ6vgsc6veJhYRVo7
hbEcy2QFGsdEq7SYf7qtcX12SecERBQeRzuUZ5KfSlrarlHZ5CDHgi41FF0rpPeE0AKCUwrIWshQ
/Bdj27AD0xOkRcZeczVsXlzmnSnuJMU2G3V2yRnzgzScac/YmDNGHiorEpLTiFJ99Z0KFqcO3ZOn
hCCebZ0lzVOyndVXs52brV+hYy+AWcz/BUMVGD/nBLIE1Sn6ILH/9UuEsPVTSO8C6ekLKGumdp0+
pEhriOP1FKcBxOm50+hXdTwotauS1XvEaMqJrQmRZwE581GuiiFTjv8ul+MEpTWi6/1XdWGdEUt8
vAs1VzvISrud0zNR+I0DbsqeXTxEwLyAN0y6GG3gnrfmsyFVa1+lW8pmeRVt76NYZlEpoyGzb1Mf
8iP0hjIWFqln/znfC6dscIiAiVSv6u8pQfE+SQSACZ1OUoQlMm8AInKTo19sEjva/BaflCbFCs0k
T9P5riTWVGJ7kVHAM5n5a6T3jjWowzoYPdSr5dpWq2h/Jo3ay28gsTM987uoLiI6CbzAR5X/ulnj
LoiH5T4J7VA/R2mCh2UA+TkCOo4htqnOzvBZJZ05dDeqEoTfrmyaAojsXhgHuwfHvj3HpI/TPeNa
fuC+SBJcZIlEJKZ9ZTAmhaX4Gyt3r/lN9sgfL7UHyLqmJTOVqFOyvfyz5D10PnzRfH8DWz1pMYhH
fxYJS7XfP50YqEi9+KdY1UCn+4uJli1w2jEBbPGWW+vMZu9uvszpDblRCwhkxfuSb5SyxaMd5gk2
7TBqU+1dRvuWefWCmCne4oQv6GsuWKvGtkkydx2SaNK6P1ZWYmMm7C1yQAYQ2V19Zu8YnYzpZ1A1
G+T6ehfwlVn+amcJy+Mk7MsJqXLXMUyKZk62hCZkEWDN5+4OJjW5rCtG0rqf1DR9yBGUjlhviTaK
jPBWGg3kMNvH0PxeINnxNHnFPP4r8hF6+zpXm7csYX/sxpPu/8DLiixQTZOmioK4OHKrvhEuVUBq
RwImryYbluePOvF2F3hOdd0WSld1oM49If5xzkgvWgljrCzlBO3buYt0WWGhYI9gpGK9sSt8JAG/
dVjkcEgSYB35A31Pfs+8Q/vyXVGA4oF6AEH5+zBwAcu+hiTwY2b8QZWj788tpdbosAiy1BY/34PS
sOS/R0rIVchL2FhpcreE9VpNOn4+/qvUxyghJtkzF5E7b52xjtGhyeSsENt0KBqcVS38Zo8dnQq4
z8erbVB1PgkYa1lU/G9vwCb6du17nU+/BIR4TmMcbDwVbLPDsGIfH3kPMVD/jSL3ZJKKjcPD3ClL
VF9k4/Y0nb1e/NMb5azKsATjr0Py1wzjx3VetnFa/Z9T1f/RSzAIgSx2eCmHZ+zVPH7748muOmyT
NmWg0vAJYT8+cTmq+isJPpOb8BxFrqhOWnYXduJ7lmfPaqg3wHS3JflQcmkgioTf6iIDRu57GfyH
2E0npn1d8FXn1v4W961LQK6o/nxJiDns/OAaAL54RN77X8IMbCXV6MVmsoE3iLnWV1lozT3MQAWf
GTyOvETvXcMxgkCXDcDZd2lCEiR9P6k38iTcc7oCq7QayJ1/Eg9UJFre+SOUxjG0UEWxhmFGNhcX
xTqNIqYO3LKerVj96CWrhlIusuEML2XwayagpAEOwLritqN/bKkW+NSt39TJz2i//11WXwxjKART
dRnW7EZcyqATmvMgnX1qbOaWDxTVM2nEAux9sKsCtvtoTi8I8KD6Zy+RElBSOaN9kdXgNuXH2uYc
PD3TW9eVafJJo1fmxRPNj8FdZJyLE0Gqpso3dvsJ7BYdnQh1bXNBuUJQHEkGQySu5NuBcSp2CCby
hAhe84R6ebInwfY8aotQ5LC01wS1Bt+heR/GoELjIcHPbBKUxQYICFLe/gzVNCQtxOWo+u/NzcjV
WBs304VeOx10U2O79VzirHCcRmUKkEZbCfgDcvOI0PR+m2MijZ3JDQXIb+LJzY3Y/SCWiDOXUzMT
KREchuXNrQc1n+Uv72EN6/zTKZFKwQONh4+3lw80PdHtdNvTKIdzVe1gGRAza+myy/sOLN7vK6Jl
aXq+lt1VejRXx1lpmQ/wxuJVX7LxkSRw1QfhpSuOO9dS23kgGzLeNex3dhnm6Ej/PR3bhXGFZmY1
npg2Vc2uM8Q4DSJG5xJUiT9cZc28GhAtSOaxi6t1xJDOOvi7W8kr6WhWNPWUiTvrbcJv/uYIVsIX
SEMOoCgbedHBl0P1+Dg5EkPcc1hxNUzpQ4J1v+P9ajAGy+wnsvUjucf0zq3mj0yM4x36VxxRDIVw
QLeQuCa40n6BcQS0NCTzP8Zly7SlBPS1NmGjP6wA20m6T+qGxc36mAb+OByJ9aRPo+tt4mwHWbmR
N0x49WsUHVBmGDVStWGr++4BRTfsmACTv8a/P5x3n5r4f4xNNvkit7P1pPwPs5N3+Q0yn2siUffP
Rr3I8gffJIWy52TK0x3iod+IXwhNdhenH6piN3E+Qf0K6axXv2GSqTXLIVPFmClHJ6ziV5EbLogl
iw7UqIcv75tsgbsf73yElDas21UTewMic5kv6bKSLT1C3KMTYuuLzuAgWO03VdgvRDnvCBlCVl31
UYXNrq59Hx0k/Pxz953FZVvOjiGgPLueWf1hMVAGb8PUYuAe+TtJAze25xwslrUrF8kVl+2Fs4N1
r9B4MERPegw1Rpkia3hLKk//8G3Mbq4KBBW/QQKmDJo/bMelbC6u6uBpuNGHldhNO8U24011Zg+i
RJxdlAey0TA1sRoK/iNIShRrHIetlheYtkn5ubvPdkGdcl6MK23Axc236rJi0Ds7aKlpeW3WAZJ9
5u0p6h2tyEPVv0e36AC7dEhYeEips9R0uBvxQo80gapeH+TlR1hvqeNMLZFjYyHStke62jtAoMfa
YiVKc4G/J6BuxOQJNqYXEhSX+JaUbCRwCgvah/cjHiD9CaMeEl+NJT5nDGGk7rdllzlZ7ai2Svw9
b1tAv2Xo591IpK2GNa1mDhvR9cnFY81XnROpIo8BBrCzNhVjVYBLF/m0Umg+FeR2tbaHHCZ4k8sx
KiRnmNCuzjk8ziV/qr6Bfh7rj6VVllEo804YlnKe+VyKvQ2KGcrmjYr+WlO+oTJjlXSD0ECqSeHL
mMHonVTm5EUqkkuwFEoQQ111kJqdiR8WC0U36E5deYpGSc+v7l6e3fhu60DmX9QBU5Q3v8wBDu8C
ULFskJ4zuJ9zn++QSS8BiJv9Dtml9ucE/JkVD+KbkrjuSKcvnAm05LyZuqH0nwUlFZZcdfC/Bp4v
Rl55zS3N8uL0rCCLNRB5iGxPk3ayZiuVyCJzNvcMPTgw2wv7fKWhgiugpVI8JGWArByQCm2B9Ynj
+YoJSVHav/nXJHJ86Rg1ospUU1S1EbqHHwshq6irKjwnGKoE1PTlUMYxfez68ecT1KRFKtZwul3Z
AKj3ObdA+f7OkxwLemAI3Jwg1IqDU49HHwTpTQ+fCSBAY5U/z1tOecLX6ymBgw0OdCS1+0RVOvEh
puW3Du+h4Eyt223bFFF10WQ/bN1M91BmoWVybzARvnoi6RUPGIaB1TojWIcNVZ9tNtDgD2jpQ8ym
Ih8EP6JVF3DAkEQkjN/YryjUg/dfrWHKORFMnlD3PNKO3MdG4kCCwozH58xEdy0sK8OrJI/PIHk9
FjcumOOBoKCbkdcCf4c8hkjR6rHzKFc59pnX7+2lxUaf/Lxp4t9UOks0HZuoDwJluOWMptDsroR5
+anmObCtOzSSjvp0bM9Sgi2uoIw8CBX0uaroMZx/7iCxYF7QGHAg9d9tr+drPs8y8bQBQ3lR2GHI
gGSsM1+h1BS987bkIyjMWzfXQsREHqZNRiTH8CN/HiG0yWCkTaMBxngpEG3RRNKowUMPH8/quLqU
FAK6E8DRAvlBL4kVbnmVjsaViIUxa8s3MzrO/8KXSet2DVFXL8ZXFNNFh6lQW/UAy9rhHn3/HMSD
9L7W/w0BrB8xL2cSQITM8qmrpTnZRbVro/AiMqV+IeUI767IvIvZxv53Ly2sUuM7IBCkwFkTktAo
ofCkttEpESJV8K2Q2TD8K/KR7B8PJgeupE6XNcqHI9cgOpDhcjKvTi6MNrsLhW2krX+ZbsO0YnSF
AmlOnK9Vg4s3lwtA21wA4wcKK+AbGNz+2hd2mOETuIwU6FzotzudpZq7t1rJaV0M9SpsiVHugjnk
ADYJsUsRAVpcd911Wm1u1OZWeQTl5J/eY5fr4Gt0wVqHSKE7WN1UgR9EkTdPuyX2yWYUTbdX8CWc
yhxgE9RgCoxLcDwyo8z73HgHKs8efIHDb2lOc/oEp2TKnPkSYC67lOSJ1eEGZ0GqiafJbtDmWUwY
s/f24XxFS72ODdSfs7EwcybPOKvxFbEErBMW5yZvqDpxF+CDd+rLyjAd5K7BqrB4HE2EP1OBRp9+
BMfHEFmbyZD0tGmKVBe/yrR2BoXiE8ZMg7ys4PKCwnZpbKHRPHHwxDMMoCrNuNt9Cl7M4ULtd/zA
olseYsYt0wAIo0eULqcQ3H+P74bXNRD0EDH2sfZGAANpRO3rP9if3WBsNg1/UBnfjxL5iJ/ev4DP
bAyGtZKtPXD4CIofDTZj/UjQO++tDl+mA6NwFvqjwEP8SW+7QWdQq5wXFNcrWO222n5+h4l/4KFB
s8yHBgHTFSkY2vBeW8X5tw7XlHYbEhy+cc+mznGJn/FolIuyC1LSl4KElr5kcHkkYRVbUrqXk5t2
WvvqU4VGGhCtY5daymt94V/Ug/v4tislvjh5N298HkEPNCuLVPRlh4aucTDTJQ9vmKEfUx5ZXtfq
JbCjOHDAceOSZp2srhBPtGll3JvG88fnpjquTVXxIMRm/lEFcMBbyykpvTvkME1vMzbR/wKRXIcZ
HrS/OoT7EVDHTeTzu4E4E5v+u7EXFlaWV3un5dtYr9WzzDKfIUzkDgF7GQmoMh38aFTkWxjqQM01
EaVIwai2b3joQy/0QoyNWXL8VQOIbOq/PddMbdKLqGOmu/5IwfZNib33gYPq/rm8P3x9LeJ/7DTp
+BGRFKGX5hqSeCbAA70+l+QTq75LrqbXktP+20Rqn2i4RgnP28biORyCt+sSQQt6mS6ycU9vmcqS
kbfxj4OdoOKZ7WKSUrHZe3DJ6J8dEbxx6kuCAhsAcXd9hy92oZPcYBW5CoFKNUVKOOk2Hb91ZNQs
da4dr/X+nAM2vCDUvAevr6V0UZ8m5dQZ/1ptsInMtkHhtLZ+ZArT3i+3PJdbsYUTk9RscV+C6T0P
0xPnHdKxAt/Xmt+NpWEQYq//L4MjT5kxsJrm4b1gqciIsoIUW4jh+c+/80Awndh8DKkHJGv7sPvU
Hrxk5rOnXnvsZLJbTTi/rsYBEPS4BPEgGplafwomWyOmQNXQ5Xo/GPnvw75SS7WLmtvYge3zus1X
zMbdGB1na7Z20Rr2nuuyQI5v0pzHQkL372Xilwk0PSAssLMIvL/KSHV0byrzYp2OZ19m/24M3Go9
p4TpCIALYAuvlHY967KPTRpZ59T1bUMdRnbErFH6f/DxSVia+IHkqFXfS0Oolok44qBwYRUmOVMm
ws1o2Mo0EgmOROu0QR4QzfvmPv8nF+F8rgmQb4mTRyrpiRYTFussDgegLzKIVucNYaJFvaydsH8S
0C2da5ocJjKp4aNwy3fQqdbF1/TCFIzDjn3mNrN5hCZbvHTjTDMzGEzGY8mRivFbabV32RZ4v5EQ
PuJl1qHDqWW2Rem8k9CZ4nwAZ8biSko6u0pdq3GMI5ZcBT5BX0C9fgETS8c9rkiSf0QI17lo2fgZ
l39mA8RE/a3ere4haPKYGBMSrPvtzEKT/6eZcVkkaa3GfWflDXqu0LOEcKdg/vGawJ/s0BZVVRMA
l4GWWAlRb731CUEHfl4/aqng5lDUKA97nU2BxI3IMRDoK1G/aVBE6/ad7UOEhMQYMFieO9gb+Wvm
K5ByA7Gx3Lasb2QoTU7owNuAvVY0dPOmCBdRRTrc3tf6TsLKE3i4AeznxhcjjSCeHX7ujuALaubE
fdlw5xAZxYacJCE3di7TDmGNipwg7Wd3ajRV/lJh9eurECj2sZacMOIXG+4jaHR1MGCi5lwskjM/
u2M/b7pGmQByyGBy+ViuGGPin3jUzRkBetYLlsieGzxHJ2n2ZxIariJhQYmir/lGHFodaxfXWXcD
271PtVXpSZ+ppYU6dwUrVLnhb/XlGyFGdBPhEeKjlJDtKBY+XtD9nGl2wFambcWKYM6iZvBC3pjw
DYtx4WhGha7tc98NvWiH5x+fegXb8ezPusWonwt0g5t5Dup2QX26NppWw06lzUinOp4vp145Hbhz
K53VktprsyMs84g0vgJcSXSKeoamFAFGesr+lZCOT0na3yyzL48j4A5exKc9IQkyEOOOadc2NmeJ
FkmF1QMf9XUCukbR1jHE67JQPl7C29DQLizpmfT/kcErJHVl35iipYg3x1foln1aKwXl8CzlHpBh
PSEaUG+puNbHlo9z9q/mMvTHMXecrd/ZYhljZtDyV5IWUl08EQiVPVUB0R35PEYg9FC9/ErnMIMG
hF7V1j7k+PHXlUHTfoupghluLPAE84NX0llPtcjWS/7QnZtJFeU5Fb7jzlsfhQExWgKSHHoceDnS
3aRl+f51IbuhfxuU3bsy4EdQilLc0CVYCMXLF91/Ix/hIVmuzMOWrK2t3+WknybZVlEHTpF3A2F0
Kw6jjz8G+cMl/TEcrVeppxNXfmHK76MIW4+juhhNk/xLAJ5uvDSya8E5D82jxKvj8sXhWQeEC/bD
PyKwIiezxvUPSEA8HPODsXPWhgm1V+GpReHLKfZx/P1vraDomuGOMFhiZrOpqFD99BmvnyKNwrRJ
8QkQE9RYTHlxYq6XJ5iz7sCunJQq92akoPRAJiK9xG4I2IhrLzLJYKuFqln/9nYTLOPlpLyHL3h2
nf+Da1AcEPmEUJNJMotlnQ8szEhjFWujSga6cFv1O4cVm/R71H5/oaAs6v/Sn7g1OGkB3XBKls9J
Gfs23dTQSAz8QEzzcr34+fqj3AcRmnwojIfX5Qj4I3K3rYmTKoZbu7i35uas/6dEgp0Fj9yxmPVj
fcBL/2YT9UCtdfWimCQUGSpUC1bbUfqiM5iCfe/CH4kcgHZf87wqiZHJTCOW4Uvo6QCFECx3SwSC
7I1Pk+dQ3j26QQB4O/PU7prDtu1BIHMQaBgzab6ZG2WVx/P0Eh7/T5W128M4HPSkcXsAlOO1WjiV
8qxdIx1JzB0ufbFSfu1hxoL8DxlcrQBUNYecFDPwOnf/rXTgW7Kmj4Yj6CBy1cHw1zu6RkN8DdA+
Xipir8F6TwAGOxFm9OLanreUQVbzjFLoXdg6PZwiBB48LQaIHI9tQajRFGKjkESihAUdv2WqWxNb
JUdGqYCz1AqeUvUaXGcnBkPBzlpy0lVO6gluNf7Fj/0iAWTHNyvSjtqqJb1/bky/jQ963lLWthvV
SGjMD0zr6+X0vX/RmkreoTfAkf3pWws3F5Cf8Mes5As8o0Bh3jr6GuNm3aAJTT9nbeYJ+5K00Jj0
pzl/C5hatofhu+e7St8Vq8HvZ489d4AqcdeB3MLYR49z+cy0oM9UVX94nkg1Phl1Oft5UdVKdpv5
kHPKcESjacNa+GloLrRhheGv13E9pQpJxoCtG1qRGMbF8LLfWv1hXIYyENsQbLZ/lVp7NcUcTrpm
n+sCSdkGfWB06FDSLsLp22cEUUHRM9CkhSuthNaZmMVNa9891CB7VJgmlzDKI8fUCn2sJwmlPZrY
b8Aj6E/ZX86Jeq+CJhBcgr1Zgn+yFKTAGNjK7NocOBmgyAzc+dv8dA5kbh/pwMDo0jda6DqXMQQC
Aou1PCRx0fbGke5nrToPqwukybwglPUcZpErAAfl3PYXGLOqcXpX2vP1llJe4A+D0cotj3p4WnYK
rdvm8xMHUgk7hqZmLUTU/S0GVBxWIDdCFZ9NmmPDnpnsPSc39g12lZ5329p/armTQySXGDd9w8rH
SLa3JQSQZiK6Y251pprq5QyJ+yX0Zz7Doak7JI+KSjTCUbFFcPS2uW4r3PXvdLAjL3B/SMwtmfbm
kZw9RoqSl4yGKACqEIvZZMsoIH0/EqgKZPHiyFgyYLD795aUvy+N8lzXjKm2cktTHXA7cHj9XdC9
mdidU6NV2jghvnEBh2CdyT1lrxDwff+lEMSbcGS9uitb6F6EDEe38oJEXxM2drPi/il+25Fq8ZZv
Ah8xBFcvNiQ15pDYKHNwY/pfzq/yPjQUmbysb/tZnl93jR9mBX/qf2/7ZsfssHBa8yice0UqLTp2
K1KB8OeyC5ewOQ+meTjz/papA0QinNyMoDioc45vpkstOdQd2yGHJFryiMDeExy1FergVWleyw4z
ejxzln+wgbMTjcCowbYMhbTT+IkwxNRYnmSNnQ0VEE3XYKjt+16om6UJdXRxvWTUG1F1vXPNt4LF
YDdm8mQxcLbXSEglmO0E1FpCMMwefqMRSGvdqRbyafzQ6d1JHx9GCvxWssENBpCoFI6ORcdvu/L7
v6oc8DTEe8mitb4oPZWJrYU55BpItoLqRvuZqKKNLmYWdBmPC9xzLzwodlfdMQd4B4/5coK+IGpW
/ae1NIE9Ali0m5GGUmq0J+uoZZwXkeUIfDlvmJTgH79lH4DMZtAiYL5nKkGWt/ecRNr3TMbKeT0y
BmqH4zHRax9LXtS0rTwwGHj1hq5f4VAuV0OlBHr8LwGs/3HJt4mTQnX+cARUIrEToMPKn2kxUZNJ
Cu4ox02Fx5CtInPzS+x6cotJYuHXoLz4tHaUoYZ2N5tYIH72BIUN+I++3FvxjsP01YiMq46auLv+
MSFxWR4x6dgtLWrM0L0aMUWy9hGoFtNWLLBiPkZ9kGG7yFBnZlrsOeqq5d5AVEYBSpqW52sT4NxY
rujE1Z/o5iU9QhCmqbv5VU+Zw9kyBRHI94n2mAg4GX2OSv5YjPUoq0dM7SAq56n2mZPVWaLg2OOj
ePaaWogTx3CfI/w8Au87VKSUWOU5Kg6A8MDodgMV8M3q1OaZKusHo0wk+G+HjTxQMv2jpduPZKDi
oGomxpjoxZk3UkVD94JQZwDwLEaTwBSaygf9GGv2eh7hjHZgWhQ/7dkbqVHGbhOsvfy7Yr7Uu/cU
MgBy6z76Y6Np72MfQx+j9LZYFuSBgbQ//LIolrqbvOzVC5lPSeeRRY/bHLIrSQm/mtBXNh4XHeXt
wyifP/P1XAaHcpDFUwPVvfurOhTs29mIKC6pnCzg5q2HycfT/j/W2h81+SCZwa72Qs009bqqjXft
uKk+vZpsJ/9Sll+qfBTqYfOMrYMjeDUeNKzUInTrO+DiKs9YFdjmg0GZKHKf9sJScHJlDgyMTNOA
H6jg1bEQAVDNQdNPYCuJI8vG1D11MkkbL3t12qipjYvUfmgo7vUsHxt4XhtMmYLW5MQf4+0KF8vK
WsMnLHs27XLI+ZCGTW6GZHgngvFYsbzq28nJw95TaDezQaTHzCrCJZf3J2zFOuheqDRzvtqFCuo5
y1i4oZ7UkRnIGIxYKWBG3a5u0RCe1L5YbjHyBR1wR4BFkue5LePy5GmqXp5fVBXr43PTZ5IEawmK
9NycJlfbX49aZ5GW64yoODYY7dXcoxzZrOzcBqx6WVUIDQyJcg3JEEQMsAG9sJiPDb4znIUulUa5
pfS2lv7NjwpKcGikULUO1dCsKtHUxx1KpuKrqAy/o5P8GqEd9xMxgN48J8HPoXTKL+eR6yXrmOhI
1zWrmGPe7er5x/Y6I44IRzCxOWJouDPloD6FsqdSWcloyxh3zuCIuJ8L2bZa1Y+bvuUZxUc3ubLb
c6C4iJNO/c+XTZFCbLve4QoE7x+wZRmJKasxovAPCbgL4VtfaVE0mWXthB9vzmcfqiv/jG9GVCXd
YonpsJxYmVxeK/saFeWG0rihIDUTm140b41j7on3yeIbIqU7xGuCrI2lxsTmfiG22rNjE1PAxnLT
wXGkJvC7RWBXVzN0ZqBc1qftcN4zUdoiS2VVYHu+bcxlqcELdr2wsos6bnHEWCspiI9JhcFeh1Oj
3nZPdLo8gCjoehsg+BDAAJ5pH7QNkJjxAzOGburLknbaY8UQGXlaMnjoY3++tyhDBqAe3HQXvurh
C8DZQp0v6gcSbkW21v6x4dy4X5VpXIcv8hJB9SfsOYjRVZoPF/hfkGUaQVyw+m9BDqFch6Qp1Oig
Xb2N6xqLHaoe4hrgntcHrtBUOZWRpYOgwd/fcIr8kFdsGKMxsOQ70E9vjzRPsVczygI/T5/UIrQg
UUxAXXL36Wt8QDCW4pCS08fRCHKEZqbU+k7R4zjP1PY6zNJ49I4E/QldENXBYrrmGLtdIjAnK2r4
58PAGzl7RD+wpm0WI7R7OFEM6Aoql4rLcRy1orXY22VN5yTZVhYhIIcvuW0ZCQziXzXg1mEs2EBZ
S6YImt+fMEfeR1ClML2u8O604/anXMIzA8G7dSi4se5W+LTUPEu564PqvKq95hNbF9dCXe0skOPx
3w6Z5hxv1WcbyX/8qfSWxBZ3pc6ASBWQgvWBapdhVzACeYRtDifoArE+1lLCGBPRfDyKpooNLsGL
nVJu1lY7sVonRgSj7Qj4LjPofm26igxXv5tDAZPF5FSB3eO7mUzffPeXPyPCmEBmrKvvKwf68zHE
cIcBfGBjCtmSgKf1Hv1ZmUIin7IxRnwRjQcpU/w9a0QcyZu5ymowS/0RPKyeF31/H6bhHc4emlhy
A6eKc/h+nvmffNG6ROteJ5f6pp7GZGDeA522EfcqbEu/CHJNocVJVctECJQn2qHcIidvJbuRwaju
97w7ZOCDPZ2EoBb7YRReFv5CT106vqiqg6QuoBBvN7NNc4CJ7HLA0eTN6cl9Bd04amlFYI5O63jt
HRVAH8prtCwxkqtb3C3UUuPWxJNbRQ0LJOiBneC9kFSZIesRaOCjvO1O1Asw16iO5nUaNUKNPN8f
ZZdbTHe2fHHNYP/dfRHam2JST4hE3Z1gCLJUvm5Yw+uXLIC5OIFt+PGzCDKi/QA/bUmNnecblkrF
FqgtCIT2KOtPPev5WgSG5fJqa9C4hPfH2xBgLN+PLDmzXjBPTZRRUFWQWdkvDuKGD0UHm7JBYKhw
i3QmHvXlEX50zGwOYviLxHCdrdAUK9wOCBINVVi3jmEs3zc5M4AaI1teKwcOAUNELSnao8zRre4/
8z60cqUnJF4DlP4ibLMXuLs5w4KNdVkz+oGrc0NuS++e8hu7d7F2sPUQw0hZlYw87py/qm+ZNdt+
SCoRhQN26jWXTX686gJkud8Yj6ou1g2AdrOEvdlH9LpzULJ7LNPUNJa/uIdA+iajs36WK3LCCKrN
ZCBETSb8ASm8kZfnmOIqeyWzVRP4bIKjpHcRNn2af/TbZgP/gl7toD/vXHl2D8oZaZs9ILNzpiuD
qlvCaiV2u+oJz3sV0tq3fuj2RVKufsFsoot0wkJcq5pvR/CZ48sQaZ+zJ/Pyx9GPE5h6gkj6yQ2l
+HQ8a5KPL0ZDnBlMBOsbPuFggHVbs0Zf/Lnq7stKkqkjiuJi2qEIRobpDfrIr3WOIaLnRY4D0tsr
roBINNMUWWWjsufR/pup96SEzSZmbaMgZZrlXS4aGd4EaV0G6OcMdGZ+wtBdXmJX9ll9oh1p8KSG
lRzBNOcXCAhjks19703WW4Go+DGELndVTR/iL+A1vtf6G+gV92J+Rksfsn9ootM6otSxevr1lGel
12N5eKOhvjDCY+rDilRSWOxw5TU/t40+lTvVOolsr3m/XhlfThzUjVoYnuPbwSgobc20qqgFzGNm
TLc0le8jZZqn3li5yxsXIBztj3eGxkMltpLSgb87DOug/6ePkDweFpuaCwHcPA81UCMPAbZpFUPo
lN2z/UGm1Pz70CcM9vt0Sl1PVsqMzLZ5f1pxS4KJh17UmdPbOefynGlF6dnykWMraoMbGtA+7HdR
ceZB0E0LbhLoEMkLkLX7QvtLbvNNcyJoqZz6Rre9JP+0WTo+9sDThPdOGTR2Jo22VkGz4ZwL6COT
/iE3CMAfluWPGw+1mc06dXtAV6v5O9fSmZRXECcrxbTWH1/u2WI+/mIqrTJsHXgJNCELWV/zw4hN
OBsLdkBp91QjRx60cEXGKtUrCHZy5CnTlfBMUFKaipEuGzDrE1EU7WO+bruVO0xyiY8y5Fq+LstO
wF6b8vjmL/xsTb7x43s49+gUe2B+PsN1nCAdJIto6ueGxcdh1MMo5Cgtol3XVspxh3+25nWCofTT
2TX8ipxWas7C+MUGSgW7Lr1Y89G370mHJSbqeHjlEtcU33+77ZhLvfnx3wj5vl7Fmgw2LndDesZP
65j19O5/Sht093JWnP8u4Y6U4DhBlFmVARzpI+eJKmpYEWNUkNcpPdKBFhpbOYUN8UG03BdYv+dr
VSLIHah8c5VdodOcTzkN6poL0GsovBlezSJhuMBuq4aq271evBOEH0o3cQq/Rca/DC6KAcz6RBYV
yp+IK1NzmApbw/plBTNqiECliQCGYav7GCNI6c/ckLrTavCFcTkFupkQdFZQNYZFpl9JHHAOA1Yv
xgWeMxZQ+jRHSvz9mBxtt1LWSQg8BvXF7q0Wn8lpayL5B3xDumHWlwc298IwQps1mZYYUkziG/UP
jqXRPoVLfyakt2+G/5zYkbcTaK53ogyJE4ek1361Cv7EiEnBEY6pAUA6z7WuZvCm40TXTWutKxX2
m+o6bbkAKqLAysv5r4SWre2Lrq6X7CvvbzkRB3mAwPL/TqOpicSYC9z2cTCCrYaVRHH62CtsQu6T
URRNZ1XTNHlFFUoBqCbnkRZ4BQMtQReMDFOuqrXXQB8KsBGb/nzn/lQgKNiz2L6ut5dCnr38ssFb
1l7ItmPFQ4eV0TaBFnQobMsHHSTpumc5+Zte/VsJSHawUM5JUV6d1XLWwq5mA8KjYL8s1iDAsa6n
E+mLJFqWc8Xh1r///+lvIfrU3j1mQyxgiPYPtpxlgmEVMmq5FnXFacUwAlZcDQLKCizXxdQRiBYl
fNxbcymdBeIHd/NvsQnIaGInqYCtqAX+0+FXipB4NIOodMnMmp3w4rTBHSkOhaoypul6MQkRtugU
dECdDinKXLc51ri778O3wtG7JCgTpvxHT6lPK4jEpEeMB7wq3kIQCu4M4ntCjgBKE234xjJYFlii
Bi9kDUNOsozWD0YW2c7N2JqewkDY0zdmZPG+QPBxhtQu9I9dp3EeR9bvqDA7gxiTwEG5IyEXAWCU
vD3K2isJoSwcZsWDn2uaHCXZU6KD/1Cg1ARmwue+Cxg5UyM4kB3063x7YTg5p8W48qY1g5K/qEqK
pWGHQV83xNhKaGKo58P5HQvXJkEPr6CAQzJK6nw0u+d1KwWcO5napjqqQzgBNb7XGHUYPH7rmzYb
OocsPY+5GUZBFVv3sNH/VBl5kC/oiGbFpb+UvrVxGEAFOWYGz7b+aBUCrMcmMwfmcZnCvDSrYRLQ
V0L7nmSRyDubnAVe8ryRRy1V3Ut4YBavTFFgqtjZjYVWVLrkhi+P5CHGFgWTIsOsHCOnuje+mDqD
k+vwwKHPmlMsuT1FJb1HPduqnrqoXKor+Pi6DFEN2DIAuOKxyYX/K09IUHgllfv7DuErMWy2eZcj
GFbqWkfw239Wx7PBAiSaG9DBcmoaGvzg6cuU+zBGsYjVAeUwRwY63OBGuLYy6Hivs/K3sOHQD5wH
5oum+fBzZKVs2HCFPXAqosYZILxcZBH/d8+2FfVMhleAGBbNkBvcXkgUOGwoRjrZ45UlVFKAnv21
IL6iIM1lqYxw0yr8rrK7RT6PHaH6W4qBOY0JwIZuFoWCHdZZQTcIisfWVx1/qJ2Ed8ZKbVQ2JhKV
eMVKPKwz3y0dc4/pLrfOfKnAEeArKhQfKx4k/ojtGcdWbkCEWmbutx2Y60tvnRJZUiqQAeqFIqc8
NsKbJO6A4INbTG0XYk7SCEmj60HE76bFy1LvdOYmFSmrL52QhkJqQCwKSTWu9R8zrVi52go0NKbn
XkZONvSN1w/q6GZJ1dMPC/PAXvURieeKw/goUKQ4xgl0WiJ/xwFeWQNZhHFTmcHS6d/jsIbsDlyJ
btL2xnxWbT17TM3coOMlByRgUTa7VkM1V2wmQZsmfFdRdo9Wi1HHt/3WluxILVISraTjSxmM7vZS
5mETe0gqwR0mm7VrkHH9cIKKkVPVMYjgaU8qKKjhC77JmfO2xAhmbAGta9gf2hXlWeQQpBvjTzNs
X7lJfafNHoEhyJg5uj/28SBfFggeVYqj9H/f1qoQRnLWI4iVR/Qmrwjod4dGJqOSY1dqyqwPy2bl
zpA4KK5xoqPsKLlti/FBvY595z/yrGDzUR//dXdkCRbjnUjUsxBpOhH3wrU+4ZGmXNUNgPsm9aST
14Wylm8aJhswkC6fmS54MwOjj/+o3s8qmU7UosJHjQ1qcL+cT/i7mVXQsMBSSTeZHtqE3JInLc1m
71yy3t4hoV82z0z44ZFtcHQHn5/PApz4vIuMprf5ZpWl55DUAcuyJ5PBSH+g95o4rFXUJiWSuyo4
0PArpq43BFKCNOsWcvyl+4dspFEWjinxJFs986A3wd0YfNY8H7yo81d51eqllww1+b1Czax7LJKt
dtUaA7THXwlI+aN6q6JIFOwo5DKirIicw3ZVm4LoJCk4Z8EClIcGVmGE/JLvfoQmHtjrKiBWXJdY
BOvkhjG7JnMn9UoqUt59QVJkEQfOvhohyGQko4Rc786gA8znSi8t4+1NFfBw+su+c0WscgZXqh98
1I3PXGdQXEcRDu0VoOLSl3Q87tBYhPBZ6FPC9kaWOo07Hl30IqKKB8aQld0RdGk7HqNH8DGAFfVQ
LxKOuKjFtBa3UTLSWDhzeWc59DLvjgXQj4MWMu5TSN0rOVR/d6HTT/hWaJU+fPJylImajAx20SN+
+Kzeu+/OLzJsrp9+W3JfQJFY2eMuZ7S2OADF0a/OM9x/T32LclQLrRWYlg6GWl09EHyDD7EDUhZL
hOoDejpWiKEq61LEpDfPVF8pUBkbEUbbkJ4wfuMh27HyNgLZMGtlpTu+QW1lO6D5+MdJQakDW+sE
lymHH9wRkWDXXLdvyuLXQiBSnoeTU88C0L73eLwB4JOx1r8MENpCJEhrKmEahRnoaDhScQUOf7o6
/R4ZQiD6O11GZvEO7mDxk9JbYoVXdUuGICwMvrxSlBLvifXFRLWLcsPlNAav/+wTkjAuRTFaIAJ9
uKFUImXT0IsCi9G3CDTEcaQpP3GbqyyvxY5s8bqzdbZaX34E2a2VrxU6Dl8ZQd1nLQj+zSyu/loi
2KcF5gBReqJheyXbqMfixmd8yOeVH7n2uY4qh22DCbrZD45h36T3qZt0vln1cfTHA723HL1noTQV
7NIh7HuXSQXjGSfKD2+4x/AFA95ofwJPmxr85tFq73/U66+5dqXnJKvGJkWslDj9YWp9UBz/Mnlc
IXoucvDIAs/N3ZlWTqSSMVLXonwLkOlYWXCLfJTOsPW0sIpt6vyfF9RLk6TEGssAlOWoxF86NIlC
mTDfZgQe7q/MBpD8xKzvkOTiLSlH6eZrq5n4j8+Z/9z+OSXMYt3i7kkGq8BX+QGzvJvPfq84F924
7+xloZHSHKJ9fz04dmTmSRr6dmpEUfT7LL76Gm3ITp9Vw3dDkM0GC0YyZnNUBhfFcaAvpLX3uO7a
2XPo5Va0M2360Is4KgzwxovEgnvgTMlgvuN654vZMmlS4K2HbRNTUYgTtM2tVBl0RsRZMV9WcQL1
svaxKIl6SlB4D1/ExDJUAgxJix5Tyw4Es2z3gQBcDh2o3UEcU9s7Bvy4JDR1MPlFaKmJnE/4n1t8
yaatBkLupZk1qZzk9NYYhMKrxbwu/AtAIUYwL06q5TN4k0CmJb6+4ZebKd9YrnU/ImiUH1duf+g9
AU2WmvTuWytIVTdl60LCaSI3cz+cDd1o0R8zprOTiadPWpzL6gAdsFRW6gct1hwkScgCe+VqO10i
v5X5+AzkdEnJJGp8Ft1cKQ3/ADdCP7KZEMUZyucSWRRa31CpWpHLXe14gye8hUhUAZlO90JBAR3Z
ngwoqgxpRRb64JmdzqjNDH1AvABeIxrcrG13yFJdOLwGJoY8LyeqM6bFtR4L41O0XLG7oQytNrIS
hZi7OJf5a0BXwdQ1UkFS+me5or+s05KCaoqeb5M07KCVjTABwI+J5ec0y/fKvteQj4o/AelMm153
VSfaH/1LAUr/pEWMuG1arzgleUTKIb8WXMucN2ewrs/felzCmRk9VqJr0k304OkILuleSTYz2qVe
gFrpAPCwe/83sJJ9+j7wjFr46tysarM3nic6FX3VGFgyNHxNAX22QzNRM32GmW4vj6I/EwX89XMu
NhVWQ7yeV1ThlLVEbN6QjK6XEyrSSZe9RIS9law7BP02QDvUxcVUNCnraAq0q+ZiMOs6V67yXiIK
2Mk0NzINjKU07WvBHzB2aenA+JSlokc5rBqGwOUCJuBhsTATwCh5DZB7gXxnTqJXqnJ2VqaU1CNg
j1BRrJA8pMS96D8Oyk2Olt6o8BdeIGvDpt2q7rxsD3sSFjT0rIULSqakICNiucatHs4eAYpnEheA
M7T5jgkQu/mwZIptfJJvrdjzFnFmJuhsjyV6Iw8uYJHAw8WdovlD2D0CY9F08pkGMa75AQXmnQvV
mBz0bao7h8KI8CpqnAIY/n1QF+qNhKA1nLlgirygIEso4iaAXfLDCDVMzvpyC38kND0kRkBm9ENA
olaILXM5Mz5V4HXdNq0+QfmtTCLiKuso1s+Hth+K2m7fae9bioqEDenoK6bkR5eoB8E8JnuzWXh+
EQxTr1LUH/9HKmHu/AB2JbkMVzhYtg7sj9tDbuC4t4joYYKKbaITVJLjE5dB1Cbnu0mPradmwl/N
3oVecYQL7V+BygPc0RkUA0T9P8O3wunnvpcC0LFA6gVAt1zLAPDKTfjjJO6+SmpTEE4+OdwrFrQq
wRbMICEU9b6de/6LV17yfiRDK2ugREVNqoRQGJfgIRf9EUZAU/j9HMvAIauCRzaAuDMTTuY8auq1
aBQqWLkwiqLp7wyCeukeV9119U5+t51xxte2t3f6h1qHItGrRqYtkaK25TuY5UlXO45dDAK/k4QA
2OviGHQpRgvOmmdTQsaur3Vt0mriIM8SMnptGHFxk2Rmcb7P4UAMv0yOjJn523ZzFc0zr+cufW3B
yLzi+dCnwOCmfusngq3OkXi+PyQZVlAzoDeKFFJWayyqPFiX8T081MWVT1qa64DJxjxIGsU8glbb
WU0Ac+pGUunguMRp+dqGM8OW82SbvO3vTBj5aM3bTFoUdbjtmhHXsh6oti+yNA3lCC/ZLS6PH2uN
/LzjwPaUE9jQZS0tmmyBW3sd2H7UVdMeZu+UY5x7BJSuZu+RmogVl8QlJUUtSPZm6QYGK0etyDko
Z/m6VOnpCFzINQWEfaI1P7G+7rBYwMAisbAtATZGZJnAYzGSoGpqlg68lDOe/Fm6uW+j7nruCdt6
kN1FOD4eL9CBmo/nTdvwk0NwqZrZfE3A9pMB1LFeldJQ33aHhWe10TRQaDc1DuK47cH4drTQp6Hk
CmNMRZayS1IcOGYZqRk6p8Bif5yEucwhzPeqhT7LYsX5Ztj/vbrvlowVUHGiFnerKidqEODgPHRU
BD91bf7Sb3Gs75VUrzNSn5gWsrs2QpFkg66uarlhYmuqHEW8fPgqww5CVbBvcXEG/AnVhoZq69fB
jCG35e6h9pj5qNL9lLL0qOv1dJO1qjQD8icKhaZGJmpNlydIg8DfWdFBuqvy1GSWMpTpq9a/48+A
vNtayz5RLLL3ke/rWfJaJifuZuOV2NgTJGvHyJmvLq4FDh5D6Ob1FgOusnef2zF38ffnxc4IGBA9
xlOL+Ngzax9N48+pZPqMnSvbtr0dfRRL7b9Yj0npc2ZESlGm3BeQC+skGqz38/Ujb+xnv+hSv8V0
UVVD0AnNfvg9VIa65dfWkaB1boNyLA9f1N7RiZz4FjrLg3JqP6D7/UgpEAlXxGFVNoQKwGbVDbWy
MyZ7SLsrQgB5QYN2wpUajYPiNZ7uLe7hZEXIItxfdH3L7SqBnyhZSK/KOMaN3mwkiMcmLShrMbJz
pnhgFU9hNA1vx4RpPB1ryXdJLfG6c6xKuZWXm5kKhskqVVeA/JVkIDylErBAbfXCV6+iLsYxspwU
vPtFeuYa2ZpWiGZd3GI9HKSlx6zFKsE2OMCxp0myTrLV66kM9IqD2PwH83vSqAW5WbBFvZjR3fPD
9gje5ZmLE8TiTG8m37DrAqePCxTZPNsBOalf0GaTT3oHJZng6Ukudlyfi/9v2NCwbMLDGaLJBmO2
msKVQYEChHoKdgITPpHUtn2SR1dW8JawD6cezMCNjlA2QdFqSxe1+Uulcs3jfrmBDhRdccagvKTL
Ie7cly8845p0F5XEytrIElW/TldltrOBYVjLs/Uv7b8zO2Wxytk+Vk//GispVGHkrvVge6CRHT/l
c4UtZYamFVtziFoX1/Hb/w8i7MX09631i22AfLzl+Wj98YDUk/cwym/D7nQ4X7ZLOkSLhEvrk5ce
a/ebaoUixvJ88e3q+3mPG1CbAduxqxiXW5ZVwm0wZ8RzbJkcZJMMc6kD5Kw71ovp2cgOzN5tpAek
ahiobNqNIQnivfhZcOIjbv/LHZ0I31DvGu1phcg1bWOmunYNgn54fY3XN0edZKVyMRd7gyiHMdyQ
HwoZwzVSSZ3uiusmhnrGbAoT2oM4A+TVjlwyRq7SyWOqrT72I6jU5vrBu0BRZ8Qh94HIkFJu1Wrm
d4DjZ+YSpBCg6VAWIf2wOIaToPiyyJqBW9ke04quMVXruSqk1h1g81et2nnbxThpyzTd/dZVYE+W
Vt3yHo86kqaOggvImvwkqHOZLvjFV726u6CTlMpVz/K9c5zaSRdRgEFn6SHOp/bQ9MVzvgoXmx+L
j/fTuiX3iLekWJBB5uu2ww8RgqABdxp8gEjK1Ivi4Nyq9jhpAZpV0IWoGcrvXv/d2OSm/xvay+3g
Vi8AfzT/QKaDd5fTxmpTQYMSGk8kN3p8c4wgt2HU1xbrVSiwLBHKOGPWul7f+2MN20/ZcnMCvWfJ
G9KyKaesLjP2+55M+YFEa1PdYUo41p9cKGPW79vjiTfzhic/O82DBogtE3az/zQHbb+76nbsAZs6
Z07NNRl1sM5X4ifO9TbMeqFt0xkqaMimqbyWfTJaS5CDVjH6O9hW2L7hW1Cjh0Q9zbT8qGSoSnOi
7OAukpp82xjZVSyP8yl7C2eUJARcnV9kv/u/+pRs4IkSBHMf674duld5mJXCvTyLiOECXjmqRlnn
YzKjDQcKJjyyrv5QBJ+1dhmCwX0pMwE0Ff6FSbUYYBxhR51lPxwHwxVQqr/+cRwxUyNjv+SHMeBA
rIwgDhFzeAklpx27D45kALrKbrF/L8Mk7N+uWr2Nbzg72H8Yvjg1S3lX5opxW3ksRP0ui9JXKatN
oqbTXH2plVdNwIeSrRRKbmDTMQOm6TIS+V0zUYfZ24mXEUIJO7iDxHyBRxyDqPr9XYnb6Z9GuKjL
JBxFaESbOgwNKqp9HxDGTSkxfkH5lQVJm8jBuMtULusNiGgALt8MyvYQVXuHafHrfn+jx1Ftq4Mb
Ou79cD2HZsQItbaFUDT99jdQAcLskuK+an2aRXafDrkrfqi3SWSOR/925c3r6YjCHc/2k5tEIF4m
7h6ikib4rjc9c6IGYLGpqOAIbP7YPHTf4SRz9+mVoimq8h7Tg0CoxsRBPPBHoumqfcILuG85iqfb
hgmdyQ/AE5hxI0aNTXFWCkx6Nx7wfZlFlUIQ1ZPtz1jH4YDj7Sxl4GN6QWBAkuHGZ0xK7sRNC0T+
sX2FSAq+C0OwpsAw+2DyVrXN4tiNUC6WlsWM7STA3LV44Wno1ZJ/+CLY6b8kmSKkBTjre5VlP+3y
HUSAJlbTzEEMh4TIPnAN0AOU4s5EnLqENGZLVGSPUdSXqTOuEGS68C3Ni4/t/m0REsLE0m0HdYH8
lhhbFuwAVyOTGJZr1xtYOJjuyapJA4m3ziZDfIhQ83uZtgG6D3VJz+BNPI2mLcK3gc1u2yFUDaz0
2+/PdF+Wlu43CfECMserhb+p8JqWNG8phj66SWjYafql8S+dC3K+Es0JZZM39+4X3lcq2EPOd0Kd
urnly9PQflIaFXmdq3aQtpT4bJ50suyH8UEZT0vRQ25MQzVhmC/W77NFgGNFui3zS7C0bQ7811as
xAFU9prY4t29cIKZCvlvKgX/z4FfQ3UaL620gtMYRpT1EH/LIHscgtRpe+ex3FOEkedFZZlse1O0
Obk1X9Fzcap3HH6712jWG5zLKnrwMwesANBJbyb8CR6isAYFODSPuJbevdNwMw/Sf31emOliSi83
CBndZMdammgRoFAKPiOdKAruEyiEPDxW2lrxZZVl7B3hg437BLbEnYmCCn0avT7U0vyJJ8x84/qg
7Fa01h/3Zq16qQAbBLlWPQ392ua2kzNuzb4cZeVhzvTp1yPMTmh4KN4Jg4+DA1rx62B++rSNlRM/
Bh83XN7R7lEJhBbZoKPnXMR5dSepnSSRSiMJCYu6UJCAUJl0Dna/H8MqXtVCSVTEBlLSS30DEVRL
ub8FSLxOdgjdQ0N6I/lEzKN1WIBV2VT314vO1MdbQKeOiKlp7nuccbDHa9NuyPnnLiEveYEbI9mJ
UEWQWE/hf1p/kSh4M/GN4n6dqeUPBgfgHdo6iakgJfp91+3wUfp8h331w46jKxNw2pevAfb/gui4
+ngCugK7NWDG33A5+H/9TOACOdgaXS6xXoGTZ3+68OwQzI9x1sSV6fpmxL19tOLxYAPlRXInofC9
Mz8oQx/58zlO3hgRegfn/oPNxBsdMjbagOazETaJpzMdbRaEnlEeBuIVPSF2yNBNk+CgLFEi51rs
5LzyqxW1sDw+KsKgKNLkQvfe7PMV7QRW3e6NY72FDe2yw2Ri9Oyf2VJ3capPHnM7ZBl++JQI9Y+t
pHUd/3JncROcu7aPBOut+rVVvbyzC7lJ0Hc3Up/gzTCEW0sfCACb9/5rXSQWjX0mNUPvsRu3gyci
QS0J5sRmp4KfqI67Cq/2TATKv8eJG4lKGWQPx8ZOhhdrX7UaZek2cqBg5b7hfCai0EcZsf9UAVzX
5ohkW3XSWnCYNugRQ3KsmgccIvhiv3ZO0hOMXfp4G4s/pV0HrEfDexeCnfV5HGiuHlCKBbtdd1tt
2Jd+45IxIhsZuNb4Y1EAGEYx+T630OPDkJ994Pl4uNa2vhlCd3rNB3MOg8MvlUed/lDOJzLVwN2T
DiERNPd8PLSlH2EN2ANrUEIXGxiH5BRJJRTovmqh1UXNNE9zjNw1np8l6RGpdLKnT49EvvbYbd9t
NHifuBwMhh/5RKsY1Oc95fXt3dX5chwHgBo7moc4xbCyppNmp9r5qNj5+4ac0yvqg2BWXGvzkDWE
lHUX/gy4lQgXbzNRZIpc/bfcekVVjAEuH5X+Zv/8aNk61By9ihP+jGCZ8nvnFVewRh53GOSSI6TF
24aHnkNRnG+oj2oRmWEV5KW3wuVwRaDCtY4PjxZv9uFqrcXme15YXTFrWfXi2k4I2eOS+V4S7Jwr
rgULX4wisei4RNvBJiO/2MyHwG2eJ2XnfWShhxtOSIdGB7VTyjfK7LnavK4xdE+/GngJujdk8J5n
bYpeQvxwP9JyLTcOa/QaqvV0YVIMLZ0kBSrIvvoDcDRg2seqngo1kKhU55cfOSjOUrwtaNEtic6V
79dehQsrdAJunlakufr4BtLkqFMiYmR3QO/cKAcG9L9J6KZRNpELxhtqmFRnioQxBDVYrZ/OVhLh
iI7M9wFv2pT3jqhf0o2WyDhhmTanYWS88xPahmvuUhothsMzP47DnjfOnPqeZFnpHL5vj/BQsgPN
ZIjQCJBdk5ql9ZziJuh4jc4caovhQJpo95duIJDwUF8kH7psE6hXCsWNZjc3dDW/603HUaTWsBd2
SajCxIP7zFkw827qahI2H1Uf3Vweqiagoo8Xf9OFbhBQn2l0kLpYPcddA3xkvAYg85nUADG9FzZt
qwU7D/DLiRLZkUogzlfRY8j9GlWlfkQuaaP2+iN2s0PJtduyymjsE9ifEko278lyDUYDqCMGC1aM
fTFzhPspmQkjgdOwkZP8cX21IL0k/1aF6qYl0gSgpbnmtUP1kooTM87A42dG2MTmpP8hDkdhBdeI
fMTqoHglIY/jcwp7wAu3T3Ml+xT1CT+hRcx8Bg0jPGil/VJXA7RKXgjN84W2Hhh+lz/cApBg9JNr
o0yloKwZ4eR1Snd3sFMT6ZAtdmq04r3tD616duKtyYAxr9SaqI/iiocuBZM58wKwIkAQdim4P03Y
3Wb2cbNVxcCttOi4n3VPXD7NQAJVJRliCMGndbeXpkfKOwPvA31SR6n5bGtKMGaRikJAtG7UBCVs
GLHMSpihoDBx8EQODsIWH426NiqNbln/t0+nQfHCip6XPK13m+d1fa23MA982raS70RNXC3vZH5W
cVYaGeSMOjgZBiRsdUbGXo3aMBQyh91HslGb7sl4rw5sL4HZPwvkI42rU9hA6v6PBjvAYGjmKQ1Q
eB1VL13iB5XQ1ft5hZS5cIheFgea85QgYN6EHuODDHLrVkq8OXE/Y+83Zs5WSX7FJA4p8Ml3Avb8
Z6aXkhgiikyjb+GiOdteeqSGGHcmRzqWS+UZ0StKAkgVsW4FHfDO6k5xo93TAdEIo6YrfwA+tl97
mZUfVprXwZ3sIvLC1R3URLnntb/bFT99xtfLUBxZWy5Zdcu8TnzyoEfnGmi3YTyUrvIV51NmWm0g
lj/p4xxPVGbw94Hw6n+bZur2ESjNzfZ/qsYqdceUiXkBEoVjU4eDUyskFqzv5Ly42FxlcwAVgi5O
KamuC9dNDg9i9Z6yvaYLn57L+ihgAqGAkyhhLyKITs3hpaagRjXKnYHVJKNYZKTdzEwTND+7CQNp
CfWj/Pus1G6RsS3e6wl2CA94aydszZV7710mPaqA2e8iwW6GBlLTsJMEqLvTfkSial+4uGjKzQmZ
t7sdNKzlVeEw927IqgG7YJIiaNad0X2fdj0BafD29eeuLaDU3o4kmhn1qRT+dgcnhbT/kNVLihR+
/hKPpusUnl9NsdBjQSvmXljYZ+c1GL07ng3dx0ikmB74vWO5khIlowSKY4DgBwiWuJKScMUM8l5I
EpSTK88Zh8apbUjWdECtcj9PL0B9rg3uiFnSGwIEuh5Z67bbv2lgClVkq8Azohv/BhpHPVPe2z+p
3x9Uwq67LhrkSLyzIDYy6G/g4eQyoUVVzT4ntQhFKAX5E1B0ELyeU0lmHDz8ts37dO0CqlS2xUF9
rV0SFtcenNqgr8m71eRi2DLPABKwQHYECewWcvg8VD2kR978sK7+2I+YCHLliv/PQjeGJ8PXbGJJ
fVLki33/Tblvm/GSOwKD3lzP5sxidL2WgX966yPBp9swyTYxrqZejCQP9KwNFAYWDyhKPns+nQ87
lcNOlD7qeIP4TYNvuagVMUUf/2AKIBPDI2VZ9eVhhuFJiNjbjUEHJulrLlh1aYdt4vHinDug+Bqg
/UAPOM6c/l7bS02+z39lhZd8xMDev4qI8SfskTVDCxvMCyDFZ16buvFRQlymPptmG4PtoNOo/IbF
pIqNdSgZ9YKmOk8CcZSLdvrVsSO9fBGiRNSUWV5UGc8BlS7Kc60DSj2SC/H8/IFrrb3lWcOvozs+
J0vHVuS1vw4B7b4tVSHvtL9Kf7ti/3A0OW7Z+qg09vQTzg54+yRtJDqNtC+nixvvDZD4zNXHHk1/
167GYrCvRoZMv5OAnovNvMxHCe6rosDqnPpf7ELBmTOQ1c3wkT1h8VXFKcJfCd+kg1tKkzzfaOGb
YHf9ZGF40hb3Xd9iDLaBlVGppzW1UBrTWgLA4EbnyPEdktc6k37ydQ6TFzTxX/MUH4xUeKiaNxUv
dnHzcuAHxKQonwgtXadMrjF5eEXhOhGsZVyvgQOJDePu6N237TD8ggcKHeyVld6UB4rIeBc+iT8D
QZ9kmCAjZEUGcjgmxXLzmCRKESx1EG9fHDCuMoyTo2hTMAxKPmGEE8+/LSHcpekwxEDYW/VvaDki
XLmVz2r+ggqRd3/00b+ci4al3X1GfPiKPqhuZzdGBg4LL+CT03BF3wRVYNmDjNgaEOw95SLpl8wO
DkzfIVwBgyrycXYUM7jl9TX0pqucNMSXFjfwdwtZUaiPrGj1tT518QLDY9bGDptPazMOFScjyFhW
UkeYVHrc9f7Qn78Apc1a4knVPzLgIU2qEPgPhToSbaY7UFwTUkQvTTpUiRQcTl8CfOYFOak/Vb5p
ZaEKnTWMcYJjcvBz3LW+nd4yVUddOvO1oCiEou7s7i9CIFDf208TclfjVJYW8mvrnQXM6xTGqRUb
4+zEyWG1VbaSmR6zxfiCdQyVzL82ChYBqx5am1w5askYaPMdXZbJI2T5V1LLmYhaqYvpXWeS+xCd
9zZDDoTyY76G/c7UgasDjOS1kWzetjUGamOPRHNJoBm8nRQtQg7uKzU8Un7quZKA0FD4ijqk6oc9
RG5AvO1P8OaL1UnoyrZxSdzUgAKEILMepVxpl6tg2aJDWhT/C8ztcteplZIp0h2ReaH2BwhF5ald
xPDCSryTb3hRqy8D62/kDqUjaJQ2GjhaybvSbD1lBshLKso8zLuc+Gl4sBL6sWCv44oCofGUbEwD
QvAMfoskV04xvfk5ZvlfXv0QuzOgyrOSwCjzX6Nk1FVbe2jP41YXAdN11M4TJtZed2+yaYft8v0s
K3L1+l6t9yLv4nhX24XlVhqCfjmLT1Itjavoi6l4wPRElsDOMTQad+eXhWbi68y0Al2RXlLyLJ84
SjfdQ3lvo2l8ZURM+H9kWXa6ArhQ9M9diH4AzEWvkZ+2nhFQu+P6KAPnQuYVMmyZp1avGKoq4U6u
J54C6aCd+hR+eblFYaz2nDQOhbCcgOwItrG2e1F3CfRfGktnXwmd6hlE5voG0ZdMt+R42ZX2wCmq
sdTZO8uX2t76cSrviqFAzm9RcFTEb0sWxzi1oJxW7kJOZq5Nd1YnEXa46zj1snYk4PxrFmvQZWhd
mH0dhAvfGsT0ovzGP9R7eFDyKWH++XNOpS1Me4kN3pzOY6rfLbIdYow5EgdprfPAQE3eYqKgno5d
5ckRead+2TdGTFdovWrK6GxUOmYGc7KPLVZgqBLwOwqAsnVPPXQ1RKC6lT9f6h/QO5i4DXDrSbnn
1rfMLsOzIey/Ga5W0K6/LedE7RkMF2e9q1OXaiS3JPDCxdFwG5Y9IdzpJdn0pNIY5Y0Nbv0TBajT
lv3svcYeLYTz6FsYtWS5PJ2X9zwHTkdmr7Z4DRnnhaYz+gPbZdYti619IZ8GCsiDd4RbBJVSyRv2
aJTxazPw5euqK02+co3LaOmKNGpOZ5Bh88eVDUP06npW9T2KwGnyk2Fw9TdqnJizqwUaJmk/3VB1
7im4S9/3lhfspZBNgjlF2EscjBnn+h0VPvunVL86fM7ZhaqzFHRhHHRHWo25EArDVBz0mrKvCVWS
0v/5WIE+Y6WANuiMK7D6NJRbKiG+7SXKfHb547FNmTxN1CnNSGsI8AKy0JV8pGdInJbvyBY1n8J/
8ZROzBSSDatSU7tj7V3j7VOKvTtpnO4pQ2fGdq5ELmcwkInRUW7iK+G8FfEGOTWki5Lid/9SJmMX
NvrKqQ/52Ev9o9j9XkmLDtErhLeGq7d0Ud4gTNzauU9HiUTmOzOR4jxQo9DeuCRqhTSKG1Jyh8gY
DOt6m9gI2CRKMY4W/tc9ecjy9fQdLd5Rqc91Dq9/R6L4WUANwBuTPbLlWwHR3IbsemXXcwNBKOnM
yxI96IpAtu7lOhiudElHmLfKM4Bf+fqBTZ/cXcpzrhPtQAzUZYuN4XvsO7wpRECOOocRo+RZI+cd
v1RDmyCAhAz6siTjflNS4BJUykp+v8gWWY4zl0yDXqzdHOC2AZtVY/Pg1re3o9TfqkTywepzaIPX
R8cY0b1wgIDLaP162pxRlSPirGrZ7XKdBceojLn4RAqkGmIY/Nh7seKjC0QAoCs1bWRfMIj5oOHp
vYMwPvn34ff6BXSDqltJnGpJ99lbMEg6DPTorqo8wBSvPljr4/ySoRwjpxojDjMSMGWu2ohIiXY2
KB2saZjpT2WBna0TbeLgQsAbDOux/1IZZY6hVNWWSZ+la64cazsYhcYe04VT9EtbUbf94jysMDjc
o7SCzgg0NIA5AqYvC6aid7PMIZwju/sFefBPLlWlssb4566R+KG//aBgNK4B331AhmvQVpm90aHK
8Jv62dqkVUC2ldVKi4witecDrxc2v61qwlBA5sbNkuGuArD7H+9uVV550lJFYNKwkdVICoicpt+c
U5mQXYxI5qaq8EXPeC7inJjMg0D7/A37Uy4ixQMIVeVH07l+oRir3933ifVfRJrMgKfHDbLItVyG
3qtHle2+h+PCbRmDkxY6O+SMMtDWh7BbrzNxAVZPkmMFSI8SQymLvcfKjctNZ0hD3MBYO2T/oKPM
HRNAOtRLr50rVbuRLNzVkTIVPwTScpUsTfXVpteBuM4Fyr1octcYzT5PQrj5uMWGHg+1wefLBPja
ywmMpZlR0bF/SqvO6o7OF8WBhRaqQTGwArWtmt1OUoFzXX/xkB2O6gEwgRdvpnOWhemDNs9c/DnZ
pli5YMmmvWEr7Y/Aol6bo6Xu0t84b8U8dP+PdnHhMk630F6+XiRXRgEq91eA/8v6m3s165Ca/+xi
zBb+QLTBAYZVOG5B2YnB1E6VySWtg6fy4mw7BqRqbWrqRAetVHqeYGK1dC/wIavnhPey+8q2Qpt8
eVqybA5MF7dfA4bRoIXRKrpxGldi7rQlA734l28CHzoJ3El8Im9F3zahIhC05+/foqcMME1wkJkO
yhHmqMKHkwcjjVla1iJGKgThR1h9doKJaESQqdn6yLcKeTVk48BtNd0KXSTjDrPets4QgjI4YRJx
QGA1ViqjtQE9C1J/i+OEfVJVcnN0P5HeMIUC0I+b04C1LFhf1CbK8CSbmT27JDocDfuK9nemnPP/
oEUDLfbXydk8+cy3iqUHgdJ/xbGxc02466V5b9aL+VgRw5bBdT/vsIMZOtdl76aLc6nxTbBumycd
atSy1RhIDF2JvtHw3kuHDRuMRpVyn2u0eqXOjvRO7jGurccVaWsytdhwZiwFHuJDThhFfGPJHHWg
w5IlHHJ28p6eVBLyuO8fbzm9xA9uDM8ikXEP6nDvQaj8mI35AiUE/ufFi7uJNU2bnugN0rg7kkGl
QKB1HSZ6GDofem5ZZfozjrnnB7IxvgfY6vfBCgha+/6uzW4vYRqmcpbUXSgdJmL5jTypho1tCvn3
lSNqlodC4lhR/uxT2/7G7KuLrUDAF9OV/G/dpGFBesfse32AyZMhXr95rk3pnAP1rNc0C6fdNpzw
jfm6DALrJEH8Wh1TkpK5qC/qcOn/mv6sUVsCzSiaTOV3V80K+gqs/2al+uFfhxkHfQSWrwE4RbHf
WhVukkb2hztP9SReSayhDEk6slA+O+CbDWjzri9neZRr7jfBv/3T4dj8Ol0cBNhlSdDTTn7v0GMP
oc6MLqrHpX+YOgJeZ9CW46MrlSKzqFYjwg/MCNiqB9lk/rJ2X6IFMj/ULuya94TOtIidMlEbEbPa
k3QqvWbjyA4/8U7+hl7xaQvdTRMlJ1tSuSJLciGmZbY+3RWVMtKrIo6QV0Uut+X1rpe7ssW67X0C
jhoyEbZRQEImh4SgkIOm+gYxddi19tKT0Ht9TIcVgVVj9egjkkn2VGM54q8nZmLzV80gEH2MiCLx
+b8N/fNLTWYQtrSChfpSo4YLx5U8yb77bnJjlm8vhoxON0kkHjZV8VNM8E6VOeO4y30SXrPnQWpS
DU6EhYcNVAKKSOuPITo+Vkr2nRSGP7TuCQeaOAmouA8lq0z7oLtTV6zjz/j75PqaaXwUpUbbN2CE
BgfPKxgTqTY4e+2724bq8+uUbtMjplqyERIOkAWcbvJCcHztAqos+8CrwI8XzMjrT60HkOrVUy37
Cj9Amsb/a4RLKeAy9T3O/jhkt0dVYmrYhutr6lKK3OUF1KYH9wvz7ICUw3oD3DUs9Q1zCys+sRxp
jkRbLgK2x5y40itc/oo50ruxMys5jIgPZhonZrDCUPbm2lfHSuvEACJtH7BJEvTS41xpy1XW3STV
/CHsGHaIrawd8Wow+wtng3/UGE0kdCoVJh64V/5e7H1aEzNfSh3TGeQp+SQBHRNBtLFsVFzmZw6W
80PtVmrpAioO9TyVOQfqUnt6aTy5qTt8PtPk3CrGXIycQaT/XY8GxRogLFrF7bYUqhPEIjVVQpYu
Ez2oW6KrBZypp7O5uJcttTY3/0qpPKMxF2w94A6YkNQShgi7BmFb40kA6eUHIN4cCnC02gX4oFnW
n6kqdyUqjUNic40U6yXCUKSYaEKMdFoAHGM6Stt47svolbfZVMegFmJBoZ3qNxKoGI+/AGHrW7wO
30/XvD/MwA9uY1i+wQa3oM3j1G2EzONvRF4yWS+bE4mCCRJhEo/KDhjOkFfj/udHLJiJqGSJ0myR
q2CR8sy7mEUDTa4z/AqtYhk1CF5RIo74yxaLgLDgMBMp/q2bhzWI+xPxte72gfFUw5YFFWylMuW4
huH40LTqWCPpieRfxkTzlD4LSApNWlb3SEsaGWDG5zetNOAFCYePqY1EfuUeZVwVMx8RDS0Ktq2/
FqkI6FTTO0LkwhfSEOAjKQWbXBb2kDgjmGWNSy5XWAWLmuaXpBqFgPx8AQSw16Ayz74hUrP6dZWL
Hoty4kEG+BQRFfQxtAAuNVUyy49x3LA/IKn8uAKw9hz+gaFSKeePuO/Ksz4uG1yllYSuWfVF/Wkm
wznkXGhwwxCYJrN0hIjXBE6w9lgUDetqt6mLR5BvX4WTC48/SC+VA0lajLrPGPP5gQddqC3XdCFa
zi29kN7s9kLUtmhnIr4UsOaDkRGLvUxqunVkINhmZKd+9xYtukCwP/znzWibGR1UJx7s8OYJdVuF
SqjODSmaakNcGvSbfMsb2P3QPvUMnOuq8eTPL9my0bgaZCbw+XhFIFtNLASnbpnahGtnoYGZ8xAS
PcywA1U5dZbKrCB1DPPz2MpPLeeOVTZO7E8EjhuGj7ji5bvG1jqHdAyENTKfjNWKqKndfhBTw+BT
BLWadYS4LAMgI0asL1+1ZQXFM86ct7MqG33j9UNKpKq/lvuTVxArEuDmszgrRtjZzJ1aJLwS8ziM
99uvqbg0tS9tkyqroMAMwdk4agwNs3szO2/7fsB3MZh3eR1dzW2mSfkJ0E8amXjrwkOjC4JF1bSB
/V/RitW0zblbOR9pKSuRhIvoyI6W70s1n1g2fa9jlDzTQlt41yFXBR4FP6UKTUASpKJ4+w6G0hQJ
qlXzmZO1ecWOlbl+t9aENmgHqTBAziNfy46EqlS9jvykCzTjNOfpiCqII11pvOQt2+F4vA7WcSoI
TKe1XG5nxKj17xBwThLtrieWmxBpvHFoYaZFinbYoqyMkf7zSmnX5lI1cuDzSkElZAug6adhX0JO
BvKIsTMAfCd3BPFd9tGI6ZXO7W33gVg8jeAH0CkD1Sn3roSnnzDOS6qPAgz9hbBmG0spn/q3eSV7
WbtXIhBO0h06sfL3CagAT48wXCTIm/6cBs2pcOrE+bqA0ug/Cn7VySkk1kRQ/A7Ds27U8On9dbLt
6eslavoWaVpTUvk4nZe0LzLONJi0oDM1vSWkWjs1vuWxn5tM1BXAY52heK4/UmiaXqQIH7A3SvGC
MHNKR3Bj0TsxgvO9BgcmJJSJqqElcapqKQni2vA/9gXsxI4c/4Z5O/AJA1I6SSbVxzVZ9LZvAJeY
w5bJfKdL7eXxNBqXufLHcSsp1Ormh8YiQhwJjZWll+BzXPM3eOOH6eFcjEhmU4Hd66z9enDiUeDY
/GrruYM36RFr7zR4NxfbaXdPPp1MLnKLbudvaIEkOb5In36FHq1q6RiGoFrq5izVn9B0dtR4VyT4
Ag28r62gwWsHA38rZLZcFq88U4m+luinRr2ycI4s+BaegffKF7gKQ+t5X1koTwmRWwq3BAdrGS3C
U/jBHy4fcn+mhxuaOTAetm+AZVz04ijJRYoq0R4sOj144+AhVDX6gNTgtzVDPQqSu1HrRF1ZOK53
Wgj8DxGuwKO02A6RFkT7N+XGen3vwaYa8q3XuA3ULy5i/HM2FGzSBRe/wu3JKsb2jyNobDXbdR2Q
+k51bK9hgbmxPSiUXO4+z5t4Q11bpBZCX0RBEGP+6rsOk+aCQ/Ea4nSMwuBWdwYvqz1uEsuv6ihH
9QjOU3JNpKwbCVQD9DbIQ4jtJEHYsJ3YuF2eCi656ItE7Nk5+eufoBnIDcQdmO3UHp16iy+WngGW
u+d5C9xLHaX6TTpqvviiGEI0eIJcfs1geJ8hR/AlSUjPCT92cXf4uwTsZixsUw0u5XH7MTQ5qMtJ
TIwWtHSADJ0k/4IAwjAWcMEif4hFQFEzuO1Br3XAOMRp2K2tzIg7Yf3jRE3l6nuFHet/BmXbjRPW
o0wEtSdI+wrjRi4iBLPM9M0XresKP7cWjw0ilaTg04XGmy60TZwjMKhqB8TfKoWY+jMB2gm3fTBE
X3PZYafHs/7tMavEDv2REyQ5XhwFmDvANIcBd3+Jv8jHFHefR/EpzfMO02WqbMOy9MV5ufFS076f
EFOHgswkaJd/TTftErXgwj+v0bBpbU0Rs4IKqh1hkoGc9Jm/ZkK6+Vzp0vj7cwKsoXH6fsQjmeYi
HxX3rv7ekBW+ow9+ik+n+Atx7o1RGl/XD5VmeCdd+V1FUjllhi0E2PI87JNvbAy4KAYmZXJNSfOO
41EqezVHgg57fF9qhjJ3rwIe3zfYPsPCqmYtGXctcQgtOpJ8ZLial3hxO1zUdea613HxQ01yEyOR
XdjU51Z+6NREB/YAUUH/fEF226ZIorhv2PaPY8JDuKsUaJfVIC3+mOvhhFY3gRRv1p+diw11IIcp
T1T069p17ef4rkwrhlz74r0zLvxGot2Xns+jgtLqJ2e21AEBfo/hdFyDCo7wxmDH/gp+Q1Z4GpNs
HLNDV4qd8WwcU7+TTHokKnmj7SGz5JljhbQodBpt9BRqiappkTbTgtCe6BTO9SuDDQuXClk6p9nS
PpmLZ27pc2ONDmjDXPJTfsoyO8qEQZXh1k45OEAZ//UR5jMMe9IuCMri4VI5zADYM52UciWJ3uds
sI2ttXiScHthSLgix8QoxQXDWVETE8UtW3+xll7eJrqP4LT7Omw6ap2pwVvfcOyp7w7sDssHLedZ
b4Kq0wLVYdgCW/b0tMrGHMKTDSpigBUTKra0iOubrH+yaisGLA6zfz8uUV779pIY4dhw4uUOfDgD
aVoSkI3fdJHpwLtGmsMpJ9ihV8Mur9Iwzn6TFZ4QhzlxfQD8NJhQicNdxJJUOysCtJkQEysh42Bu
OrQstBePvPwpQVqdvFWiniWCWS7m/PgoGhcio2fKmTtF4KS425YCvwSbyKS0nemJUgSw4uSOJeK4
4RtLAlzZXU97uqpYSzUUaHz3kpcrBqDvw55ZnY86gUhVLpV2YEIgcQraoaVo7vFf89UovP/j2ZTT
uCp0zmSXHS0vxSj+6Fa7A0KtJSiPvn2gndoSJvIkqAeh3x4fj23MNbRyJhR4gAisAIdp+WPV7OZe
0kvK3MkJDBANxV2FAXa3WoSc7XqT3N94UZZQbk4pGULo+6rm4RwSzkKsgxA6rSlUo2r04DBdJcMN
1cRziPZI6N+xAZNccmZockJIrr2q4HHmTw65rHGJLVK4kxB1X79EVakvU5fzdW2qsPwPbXXSI7Ea
HPTXTHuGS6C1Y8Dz2Yu/hswnz/GLfuj8YZb2bFhERFCIfM3lv39ayZVgqghtxtRr4XLQ4WmzBIEI
wKBN9rpGLTuPp+WCoyOL5ZPXIKcOsaMru/6IWHpG6Ni/sQ4Bdwy5eD3Hratd9ddVR4ocKjNtOtj2
/OW2GZQ4FyHFKPIwV4I+5l7WwK6JKWZy1jrEm4hCN4YGrrqVfjTLZ+IZCJ3V5PfrwApAyZfAIPev
2Xy9Nnd5hMMRMRf36bg6vSLGJNKttiPG6fnAzKenql/JUWO3uLkNm8WQKBoDfvb/ceZ/KORKW0kY
/kjZwHcrxOJkMmMfNA6ngUn4PxhI5/3HpVn5xbUc+WqSCx/H5BfFwnMmob4lsBwoyJGjXG61zpAM
/bKwS8oPUSXzXR1p4U0kZB3SXRUoGhMjIx1gW/t/b0qXq5bJmusDsYd9WkPk3/iAFRL8s3z34PIl
ZxUemlws/CfYjMZiTNihfWD+/8iU8gdP3IX4g/s8Tq9Pxtzv/pgPCmYdQuIjaxEnY3/DqmRK6DKF
msARL0gjN4Ogt49yXUTjUJsvFILV1EnQYma8TQv0ryJUyHfDaIgQ+7J7rQa3WMrCsjxBr+WYkC5u
4j2jwvB8pRgtRJV4+WOWOy2vTcFwlSilhbmax3AUNzqWX8fDummMafa/1fNoAJutzTOIFOnnLmFK
ICu2N4GMyhp14/xnwLiVVYjGID3pnrXURIzIOfLa3ypcYpSKjxxBdWIi2tK2Z+nrgk6l3SirEMsg
bmnkzIhUDYmeiJDkODevbsMvcrS+i4qjCodhj5mS+4zf83uvVzPRDM7XaticfPe72YmkO0BHfll2
l2WI2aYSfxIngRMdUPbpAZHqt7Tka3kYgEfTHAmJnNBAEG3RSd/bqTWyerMqWdV6EJ5RBuTx6z6T
Eq20pCGsJ1ljHpp7jdCGD0Kj3r9gWhCBlD61lY01KuGOnU+OSsXzcEs/G43DcQRwTgyB+BddPCCZ
X4Po2r+cLRjLrxgb101RXTudEt2bJkdhNpQUuQpcQDCHwtyZ5ZbGBOGeilo3drVV/YoOkd5NvHq7
0U2Ud83GWwc3X++aSxhITZzTcH5ivfIaJ3z9z6UTC9DHLrBFKO2LcBVWetMGR54us0TvPDv9SBoF
P4ff7kBuE3J8Cizgf5wb+6G+rNCqkWAf/ERUfiLt7HQft/Z7clNe0H90cGCxn8W3hOShZnDBPiqz
buyRJOqsQrSGKDObje92YAvmD4e1jz5RZjlJ+sP3xaP21uiccYSrbZVnQdB/hkpZAFsL8RkHovnu
2FTiMwAlrgY2YHGd7GBoRYrBhDtoLBQ1bPVrLucgBD/3Z5sODfkDTbbr3/E4Tt1d5QTSWxe2K15V
vBbxv/POvjUUUJMMEhgIL4Si/6BQpP1d8SwElQYkKKgBhCExZtg3Q3a4LGvH8fyYEmSZgsC3AUhX
ehGmyIAQuI0BdzzmNC/8i/hQm+lXSB7OGBfotym60LqZLA/T3ryi7eklb0FM1ntukPLAKmLn2G/p
xg7JYKUKNKF/aANV4kAC0Zxp6EcbmzTf8r62QzqBuwu9ZrpR4q2hd4FmoHQeA8q0aFDJUw1bXyMM
b026R0mp02qbE5EsoadDQT5GZa84GiK0MuRAva1GpV3ojrJxnZRMwcBDeNSuGjS/JxgiN/x6HM24
EqVsWRN+k3tac2JERYCI4lIcPvx4A83YEW+P4a/OZZ30ArvQjWaDAftJjMQ5e/Pb2nDz71C9gJ5y
lUmV8lZxPWIsTQ1ZjV7TaTPet//pRDrhv31fkuOlgWcKXz4ozgXXG2C1+7SUrKf0Pl3SOiZacD3p
ySf68vmNLOKSYggX4pZCQkB903BBX9RKYRNpGn8cgS3dXl0ctNj03z0xKAa8uGLtqEWkbmkwQWpz
kpRHAMd+ZapyCYzuOskuwfObvkiAGnnnMv0txd6LOLh0hAqw8kR98Th8gs4IT/KgYPID8Kpb2Za/
Stin/cquMbSfYOD2xlgWHo3n2F6Oip7AGJiqiujmL9P5d7s/ltYG9CwTTAc+/bgRz4yocgRrliMU
y+WY2qYPscmyR7gkeB75yY7MIjub74gudId+sfblxss2C3TDUYA5Tocj8rfyPjip1GmitibwGzH5
sObUZeBwZYqdiMzV/3/+1rQEyFQGd3tDIEBoBsAS7SHHmXu5T1a6AX5aQgvQfhKzQNIxjQgGyAhD
od8YxdtLvchC4BGnGpWf25N32pU2QE1Tlu7MhnJgzNIRipjb2xNsPHE1ffe/tZMU42nCOFaKoGVd
uRt4ay/XxaGIc6ar/8oQkc4sAtOtIrl01koQHdWW2Yi2BFRAcwGDSBC32/R8ZpnP8iwn7MYKwIG1
XVOfLngu4y8EK517I6/udoYVPWRXB55CMUGc676uOYdywL4jFWqQE9stZuu0KbV1yOkq/pF+PF6P
ojiCFWyPq45Vj57tiAe7zHHNM/YNnJQ3/E/YEMST9W/PLMplIMWwfTBXq/QlDuTWP1Z3sjxnSR26
9zPXnGOoREmbcy/lNcxZwoRVMqRiS+OlxNqhAP7c/f0KFKICJlptR8Es0NUoPJ+yFCs1DDmtjTNQ
lwofWGjoRWbjjYrQifYwsNTrxoPA9wbv3KFun6ATdqto8b5rW6AsNdB7TItj1XYeSRoFxfkvG9Qe
m7AyjIKFXNkqywPF01zQBVmRhIFo02jERrct5c08DcuaBW0NT7fhDmqT1SGReVJlehD13/QdTuii
gwN3uyVY5R+FN9g0mt6wC0XsgsMj2pHw4ne8LA6RJ9WnAJX9thF8rgvaCMcI120DyQfiGEf53m0y
CbmR1d9FOKFD60LevRwJfegLCIzIpcpLAMldJZK1l0BmAK2hwg6g9ZZO1YKO+FbD+LLUYsZad417
eAzKMFdd1Cqje/yAlELLnffVp3MkXJG/97zIznpLZTZLPnTiSO1r1wv0soyUNw98ziXedo7YjU4q
hiVVZRA7giKeFpBXsYWN2TCn+2GF2dmXOOGZ67ivb46eRqYUXiK0FlvW0/Gv1pfs1KZUtKBgdwTP
l2rTuz3LPjoA2V/o+UYt2XluNdsCJsYfpor4FMFSf7jBMh3t3s9EoYF2zA2nCKiiRQd5B+L20qGi
XPikePZyqDEgCVUTDMdKVhX91Ig8OQ+nqhI+vOU5/pjf6Z7I1U3C5dqQDOWLSG73Q9Q8SaYvYuO/
P0u6+Zxo9jF5fF344flkUSUq/MtzyoSy1NytHpMjVdtisNZaXJUk7jxw95naR6yDXv/BEmXRcOjm
eYdFR9KMI5eWVNTJTjCWnJRWUBrnSnjN213WX+bmVyusH+y6kc1TGm2peuRJOni1XKR7iaGdgldz
y0snOuiMeW9Uzly9NaWxEdYYKQ4zeaO4VGKPZHgUC8nxnYpVikM7865asOa3Xx/H3V2gofjnX624
zijVT+ouTNjpLuAwV4UQCMYBHTyXfqX6FFRxifjksi0pRz32u6GTWfAhWg9b0Gf13gVGD+XCACE2
FLUs1+NJTaqGNjLXe24ywDVQyIWiGYmEcH5GajiXxlgTdb8pTKiTwH8FmuRIdTqIQLG0BmJWLDR3
PN6z7qW1rxx3aaXFsK3zmuczVRwzphiFjf4fXNkSPLcejt8r+hhxz/Y4kuk1U6pctlGuB6BlAN1H
sLVHISD9maljsKIYLMr8f+QwPJr3mFHPmtuBaCpIfdQoq5RlANiYlBbUIS/v7g1BwqsuFwCzJme4
pE1Y/tifiteKDkUvxWX+tn7rLHgoCxttidyKt9tPVTFMsVE4OeBDUbygjbM8QjcKcnrEqQhdvymB
Ul69LSYQawaAWI097TQXuT1u57ZIhlDNvZz8KkNGoAG7vb/faE22yWq0LiC24ap5MXm3Gc1cjkdg
dx9KtaJmPp8bnVYLldRAbC5gdrmaJy0Tk9Im9ZOdjlp9GMNetsztn61QtztOp0uzahGqC2sPg8w9
5BEkwDgE382+KY0htvjojxoslwBeLiEeKEwuXlIyP6gjw3QKPdFs80VP2FkmYcbbR2XfxySD/rGB
ETUPwOsQc1NZJY7Ou3tcCvnwS6CcR4ZYYPZcqfnZQwCFfUaUIQfEtPXBdtm/vQZbADML0sbiZC7Z
NIY8WB0R5EWyTURp7x1r1xeYz2HISAnEcckQjFakaM1REBrj0pZFnyQr8rjNCSdpYG0rfvZ0bfrb
GNEwTkwr5bb8/kf68j3sTFv4EiOOlDhtjIds9VXNWWItFZTeVJBt4i4zr4kxm1+PudcXxYptaZdo
PP8OuA2eNnCKQKi30OElciMweIy8fyEiiXKr0y4CyR0sTsCayrsz5a+tgycwbWT2hIqbxQT/4Vgk
nS7noDyESQ3sT+QbKjHnZPUTgDlG4UTgnUcqF2EPo3+fs7d36h4cG4mLp5dfeQEg1WBAK1qHVvx/
OBRxuQ0Mj54qcJJw3r9gLJBIlXEcC6xH2kpKOv8l8GSiFOlxWDNszXPAsuooTZKrUo0onOWseUWw
Zg4TGlS2kBTzy7pkPKkaUYDxDb7qFR1+1CKSSwgxmoW9MV7YDexI+qNyhF65bGlOy9MEKPG4YYmm
JUouXyfeAMoEqEPCh8wdNdmBJgkQfPg2jfdRIw/b3z/Km/1N5Qx+0YfxCaOU8o0eFGai6Qb/5Qae
hM9tM8JsmuXzOOf375Y1eGBpFScFlsJH+zNpWsyTX9XxesAQc0w2XjoNTtLVT7UjT5ze3vxuCLCj
aH8iOZrYvWdXcKqlk1zZenaGEBSJ5bm4YIQf+ypDTH3z5uPRwB0hA9xPbYp4QqHploEJW/Jrs/HH
FglOWQ+z+u+2Cia1+ZBAgBPp7ES36ZiG0gnm2T6SPDrAlD3yGqk/4FlG+jYUOTRg+9lNWIG7YixU
7z2U80kTGbSDdFFBqjSmVUQE3wVjp7VoX7tz6LoII4CGc0YmGOruKBXmm/Bd6TprlPqUDkd8tAzj
DpVB/7M0/AhC5jB5x48hUQT6YYI+f9uUc0MvOCiRyQ728+HdLMLLuE1tv6TLOio2Jjp1KIhoHFKm
EICqcXBf3ExIEjD+UWU54BJ88VYc/rATGf45mhpS+uht9iyEZVYs7a2gjZk9+9eZrNiw71svhXzO
nz0kAsunUOhnsllGeE6YXvQE4/6iiieyk8P2WUh/ORoVjcQRtiV0kUfFE14I+fDTXkuhD4waEVfF
xw9Jbgxi6Sm8ubg70QTSRCt/NGrNLR0ZQ6BIPuO/6WJBL+XMtDZ2mCXlYPpfRNumqn/Gdn0bxsI1
PBQ3MDl7SmSqcQcBBmyrx9ZcVi4aDkZTgsHOabH3Pm+RxZzXYv59zKIPM0mbTMA1C8I7E1EGY94g
B9aQXNsKzB9xUNDH03A5B88r6FrPJUSa/BGO0SgohuOxwERNsXNLtEfp0x8Df2/P544IB+VadBBR
WWM4DQIFXwPlULyZL0m14uvR8kXXjh3j3KlbkYM3Wnou3XZsTPw1c3FOHmddgxiL3YY37gh7GIMC
jTlqrmffo5+TmQUonMfG/HGe6fDsCf81wc+LNOhwrx2hS4nzv99fNYE3+k/kVOZxGfra4utq1m5c
xQOh0KvTMS+aRPOWguN0GjbmVso4UUMrmzMNbHFStgc1BcjqoCjv25+p5Fnq1wJoqPSdSi25Qs/1
X3Md3QM1xPZHR4PJv5LlzTEZa2nXt+pwAfm4kK0ZRRNl6aoQTHAd5vWUB33+Nd35HkHLUxsRObWe
+u+GU1jr02vnC1JBt3KkWNKrn6xJ4tVlffjqjEiOBFIlQuXq2XENMHQwreWY+scFRKvShYNbBRqY
4khLG0Ag9gb1lxk+PYBFS+Dc4ltvFN6KupqutPv/HvanNOnLxZtG0MCjp44iqEDfL4hy7uPgrZfg
9AwQ2LsS9goEZZD84iECT+iFkDaysCmbBpdyaQOFnicApC4dYzLHgGydP8w6uGURjUpQNYuo3tyI
k06UbWp41Cv27y82gpvvWtA+N5yx7pWJ9iReh6LQOJTt9Fr5WH5H6kUkYFJ1eEflWSg6AskZunDP
WusGLMCQZzFedrPeAeS8ycXYaG9LG0CaObaMO1jIyfp/2kiGJBfxgYaIq5n04dpDdqg90KIdt2hS
hMH38ET8UX48C1c/A1lxczV5zU1Ve4L5uii8TQ92+7zsbioGETDHtjE/e0jIRNE5DpbQ8nV2Kz/+
1D+uOa6XR66wWiVpy90wNcHxNY4fqEE2BKqs/MKqRje6yCA5M3XgTdMn5DvXevpWt7LUlgc8jBGl
tcZfHZIwcyCXXUuV+SRjN6cPuJBVSt8JV0Dfgb8mWKYWSFe4RbH9kgIntMbmrIO1Hwf/ba380n4T
6Kr8CUxse0h4BuHxxWYG4g/3QLAgn6ULMNcVEmx7kfBPrKTdBWdFYpgyvqJEw7us45WjZcHIviNS
lEbIROWQ2gVQQGiQCh7dd5ardi4PdvzFkJ7Q8qgd0cxsCAu6RUj6PSNHxUEVihr0EbttsCKaUeLM
rvPzzl8pBD/nzfmVlVdBHccJBcu5WSpdYmLR6Z0TfIwogSCNmz4Hfdbq7npKESBtcKjdfif+uw43
QLfxIjP1RJQw7xTw1ZssffiBhykDy5Oe4gX1BXs+buX9ItJgLAmGRZ48dNX6bzUt+ombt662HxLV
WMnyP7Q+oYgS4nwhO5ffmcsOaaLe99a/Q2apLVSmOwdIMZswbOsbObXbZPCGRheMehUPNy5HOabk
4hMIwaGOlqQfAdYCEawH9Cf7vslJxXyzcjznIJxgZj8Ie/KJ8gMzM0ncT+nVHr1WnLM/8EQ92Tm0
+/4zGJ29/MAOqYmrFOlsmYh6P2rinaOAocfxNMlIriY5PvkWrJtocSI1NorMNJdJwqOzawqogePB
U2L6JWkYI7b3HP8ZPOaV1dWQC0MHrcyP+8CmlrTiFj7zR7d3SSOJRR11K89UuGIpyNcH1DxhsfaD
MZ5BhvOXWnOW4ZUzBmihoe2rNGJxqcEty6v/uTSKa7Tp/zEEDc485N+eQ7+sDU4nmo9wwg73Z/xy
upZ0OczGE91dntdVaCTPUJ8vGddXEFOBYBCIuZ3tS5CstlufOeHnUkJtTy0KOTHMrBjuQjOXoXGB
mkHMnpqlgOBl8xVSKnO9cQGaCA/4/JnxUvWs3eBiO1D4H/PmDrA0TJsAm+1LIRe43nY7Cf5LhBCh
TdXfG4oiOForKLDjR0Cw/2Hsh5SrdptPzvM04PO1hY/FYYKlwEVdUb8OUd/6cYEt6x2EgIonpck3
DGPM+xIIKmPDa8kRDjKNtcVyxTBUWjenSh84OeWsHJcgqVZ+WChQcew0Z95OVmw3wm9936JDMnuJ
6ldHbGFnGLBgBoIYL5PVDxATkOUpRro5Cvyirab/JwBxiblULBZbtBKRZyxxmo8hT9rK8Mzs1YO/
BbINX5ptP2bkdhHC3G84nPd4xXOpGcAHJ45PJ0C/Sc80mlbjy02xh0V2ubNsIkckMbKSo4/Tlw93
W28pFTXhHlE4h0tWzApFQGSgYT+fwr96zksrxmxOHKoVLvEOPi9+SU4bAYbJedDvOWQ2eClMpSoE
Q1VEAta2lpHkHriXJiz321Wso2dm3vVBojl7R24nlBsdiRjkkAlI38rRtN7koDXHqo1YwwlVSf7x
RdG3/utyYorhprzM3wogeTUYMXLJPqT/T/jY46wNyzBYUIyH65WeYWOsBXrPuAlohxmaeHSXB+Ka
JPzD88i/xWsYo44MnBKe7hLQmCg1dWuu5wlMyx0GpDtSFK0jaTvap8buxkygjM3h1opNpylwBPjv
eq4+UZvkExaA0BUuBaPyrJCRaZUQzUaLetg0NG/3vWIGQBANfcN8aFjjQWS3ACzJF2KRVE23ALQI
KF3RsNGXvOR2uK7GcqT9v4PMEaj/NAJmAjQKIeBcjmRzjKTVmC3dUoFsyYOjhnnzwnDIL/5ScQw+
+xye4QTnlf9weKXm7gI1FVWiquS3xsg+p3eN+U5YIf7jylDPOwg5V1lHbLpRyw2OMUUxvrtq0obu
PzN1LMtukpg8NbzTJlNoEOZylqcq1Fau8bv9O++rdFVf7jUZFSgZE6caIzmBLCiDKkb0S3TOsUoF
M+sCE5uWkvxUnmb20JJyPK6SD2LF+zc3Y/qA5EXr8aUj9TemaDbUrgsjnRud/z7Z6hVPgHNGG/GV
1XRyMKWc841brYbKja9dB9b3ajx4x/t3Ut9qgcIh4N7O2CjVKRg3Ib62uc7IzGusrUn2cpgPeesj
Zr4qInVcFOCCIqwMsBQ6NSizVRBo14Pt0iTA6seZ5VvVZpXm53n3i+tf8RiEwHj6R/mBzk7jp817
DuYAP4XlPSm0Tqx7+uaLcvJ0IrRsOWE00WQ8Ue0dIDio6Uh8Dcom+xHMu8VUAE2S+B23LMoF4hcR
+1uzN8qgXEHM/BcLdRw2tD3kfbMmN+S31D7tnaR/A+WnB2AZjVe+XnjWyhhUGbB8RqP33YJa48hl
Zah6+Y+6B+d/jBISn9n+biAceG7f2AApf4TOySfzhiRNA5Wb+Bne8k9oSm+XiO1h2bWePaLUJhCq
89OnzAGFr4v73tAHu2PwBZG3K7PFnis1v1w2jby+TVJ1PAczHBwG0MaKEDmwxLykZcTxWSUq9dpY
8+F2qWstdKS1qsG7BqBXxKx6kp/akUxNEN8d+70cb60EhBx8XHV4FHSzR7lQC4R33HvmhX5XIeHM
+mJzzC70Ws8ycbI3xaoVnkJUExIcvZspSyncfSugtnA3acExutJb3u9apBXkT1zEeP2sipkAfFLZ
/+OuekXhHSJiipfAS9hBGITX0vQuZLD3A6+T2xXwupfLxnTjO+pbfGkrWU3T+jAUz+5Y/jbjFI3G
jo9jV4lQW2H63/WGnJ38e6rgYPGOTTzehy25HX3V1M5zmzsXQ7wpgA0OsA0gdmq/li3yjsnCTEUK
C3e8zvf6szbZBeDVBAj8r0Dq9IxNY0lAY3WjGDrpUvS3Cq+ONIvw++hYWsE0VIVHV3+0FNxeL0ca
/wY57TdI+nLCaio5bl/nTkMR4LRnQEGQGpdcqQtVg/M0+oiCQXJPY9BlNgFncJi1ZlmtfDLj0tO9
ZCk8TZwOjICkxew6FUj8+I0DuBpsxUKsON5H3wxbliGV5Ih0mba1GHpyVxWef4+PJz2BfpXoG9xD
AcsdolWKgOjyjgZjs8qWruWKs3jKVXidELYjA/NqTJmi9tNMEOJG4k/YrAFgbpTIQ5BTkJi3oOtQ
roSVtYb0O/nkPnkJ2J9nTZGFO2x1478Ck6163OhBbu+stYVTbNGZazj1+rLzANHRJMEaukkirOby
rFHoFpuN7/BXlWHXuwlpmEMK7VdhMDkVZ6RmbDLuKJm7IEzRyYqIBiVsTFK7ep42VZzoGI84Vl9W
PnWD7mBKYYgAqNOy4wAjOPD7gx6M964AYH7pq8VkXv7uhoVOMQQUiGoIhhALepsOucWrWnQNEhnD
Ol5Qok8QiXQyKywJLxWZFqkoKLdSdkbDHsM/rxDzntIznpHEyWO1JsOKVOExktDGMriaeQR/JLLK
i9CDPiKCxjtzpUkBsFAgiogMNwcy+C+yPz2bmJqtc3+1qiywluFYMGYplGlNl/T9CwUonMD5Jvu9
Dzm9Z7jAgDok1eDPa93d8FyEzCc9eDvfSy+wcjuels+POdI3OVgVDTfiZvDPyrixHJkVM1MHa0fH
OX9eW/gIOq6rkNXexTPOgBTHCRDP11ZX5KLLmElO/hZ6k9tUlMBayZBmBCw7EIXlVsrACihAN+My
AW7ojClsaixvKz0IpfyNoRIzkcGtWU2t4qBIc/xULjPIW4OtofNf3GVlOJX1fjD0S7rfv4jbWdVd
yB3dRY3EdNNfGixoCIREHzWn3gFNUM3/rOt8saFU8QVXRKkQuIWerkK5MEm3lHztnqgryKq+Akxa
Vgawc6S/qvMH54aKwR0U0IT7pSaOCGZA4wUzCY0O7M/EUNaL1Cl6794dnbFa53BVMCGwyCgFm6W7
EUqvI+FaD7SG3rZ3gsr0VIV+j2lNT41Jw0a3y88Ejc9aCrDS8k739ASbZbrIH/e//PlvbxjRfAcl
S7LQaPArqqGrpGbN1uDIpq7ai8gGPoYi/g8ZJTkRw7Xoav+NiWchyiUnt55VlzdJLaEdraiicmz1
nA0XejCAVnuY46Gg4KmwAhb9gDepNEQk2/OrnD4+2hno+orN0RQ9Kky677bjBcXkL1ogjd+LpGs6
9AdYQf4oYNwp8aWXVo9cQQHmr7wql1fh8EqYgqexj7dts7LdL6sUPyvo3u6m/ZXWR/vAytvArzHv
gFADU0PcL9CVNAlMm67mZiZf7OxFQY5troUMiA4p7M0UjriLsf7vOaq7YUyeJwezdAwvrfJqijKY
aGx548QAChxtPOFW8hpXfZNQO0/S14gyHMV5A3TS608v3rZKmu/qJIJHM/dNSBLC7jmS5ZZr+ytw
r/Qqyv8e52gerR6BG+9Q42RAe5cI6+H+VtDdc4e2Vnoq12WWom7DYRN9iMnY7symIxnuHOFaJcEW
A7VpnMrNc/yoI6/j1n751tX9Fbau6Nhl/trER+Fnz6p+65YJaImrjKtWac/L/jWmrPe09d6dJ9Bd
33i+qQsb1qw5XW5VU/4X/Puomz/Ip9xJThE4lil13gEpFOB9Kmje5TgHajUDhTkDAAO36WK3oSCc
GmKfLDSFrCuTCKurYDDNVVTARsRP7lfIyTrBihbG3yHBY9n7hFmDZlV6nIyptUO6NPbJA774ffwf
3EG1fzrLhMbRgFHq4jp/2elrXh11xXppkm8OCvlUaelK6SAqUqLqoDZuxdwZvr2NeAzYDJo6dmxa
aRSZg1jfG3vxMPJfobfGpZmIsxOBtVplLNzM2fSm7WyfWiGTFejNZoGzONIMyDdE3p1lUf8xPo/j
NQbckLlTNlhBiNdimblooI3zS7Q7jopde8kL5qC0PzRkPCKThhHRA5LWYwmqgbJpe7wJyNMuBihx
CTDFjUUO848HFKiYH1dOru1q5xAnDmrhYzLlZketNMQAquVERaB7IbJkf05zH+v9nwSNpFTC/6Rk
SonX7l0brDIozn+9oGdvZBdVJGh8P4J2cNzMt3hxL7hFmOuZBqBEvogy8cWtXAh68x/otGf8tI8c
0O85cF9g0zJl3mMSYUI1Mc90GKVLvu9d71wT597+4w4srSAJRPeE2AckDETNyXwxZ592n0XlwoGa
lt0FpoZE33a5baS+6CfRr6A2g2MU01JmjCrUQFH6MK2bNzbNuUjJ61ycQ+p5wIpD1WzylghknIqy
WMn/CGaCMnACG+RAct/KPaHO+LkACahkXb87xFhI4aIN74BBbS6IU7q8Yl8HrV1yStRGEamF2uWK
PT23cKQssbXicXnlw0oKtErbkSO7ylMpa67ZVh8qIgwxDRAtsY8BsTiTEd4jIoONlVhxhyjXbz7u
Buavm6xeh2xnFW7BoE7Xhr0/nKeeAXKLjkVPQbNCSOA2UM7Ae6U+OMx4rhjHaA8/ZPmz/GUImesi
KLRQ1Fre0lb2SqfEIc4YmF3uAmBmmNvI0kDaJLtrluI52I14T9lZMnOHlrXXELV1bl0IRIJVAw/s
KpK/yDmPN0FPNWemDL7rPKBXkdlgLAqUczs4uyT1TW1q7HKwfCtQYec+0IMuB3yuDeHQwDE0Ig6Y
sWa1D/iFKFbigkIvjvX1Gwb4adUrfyIMFke5Au+SWEynS5K2HeZWnpNfl4sujRnxKDavAfLsuOVl
OUCEkyZkoSkoYphYMPFQMD5aYfm/9Yfr1qBFRobJWX0Utr0qt121AMLZyE6elFLJ7yNuIgaOtx0b
hJJ31GetwExrR2cF8Dpv4g7CbTgQLyFIyrz28FG8D2V+97w89WpqH4nvXaaR+MkKMY5l7WnPsE7U
kVDIUHig5R8YwG4PtEk4su6atzU7gYNINbhXR49R/8E2rTrfg2FKh7ftlcNkze6aNNrKktYWw4uX
IhZ7aBWkSZcROQsUS2vGxoAYKm7rFPBBrBQbg94mtHdR8xlYE6tBLvyLtKTp4wvkSA/9vuiWoOY1
ZBwMo2skq8zxjMk4duuLM30IXWcfr5KhNd0u0bAWhpulcJX15MfSvDnaCCQcQ7r7Wm/yuMEEPwT0
rKSriiqvfIe6vbUwiD2KMrbAbuY5O7HFFFStRa++tlFeirXFAJjlrtdTn+eWD25e+H+mPdyqxogS
B3W2V1b7/OEoJj7G5pm8Zh6fgZSVd4+3RDx5CnBwE09b/4zwbHyASm01Dg2zeq/9EPTq5IrkgZnP
OqSI94HZ2Nxq1ooYwjGtvKDfzq42rRWU0QM0mPoAnU8aWzqFINLJ4LEut/VHpNpMlZZXh7skmqXm
0GFqq2MxYfFAGvWdW1fF/naJ5oWhOo5XWcEML2zWP1oE+qsZInPAd0hzhe9gklEMGW+S/90KD0DJ
TYcMcAwfdMK4l86OyBqOR8ZXNuDP+ivFx1QLxJtkwJTVflX5ZjWBqyJ4QZfztX3tQhyfdlsOODGk
HK12rfIj4uxTRuZP0iJ4x+Az8A4v9BTN5ZJBcitxQnZT95utPw4pLqxA3CVd17ZbL33RP77HsdnQ
5YJWuUlNKyKJZUgdZ4mhVtgEN5JRvKU0R2HPuOghnokr2flFjSdexqxwPsHoMKQWGCCWyC7+z8ef
JEfsfl6s+tD7IFU56QwmfPd7g9voIGJ13lIvEztPYI7z3emJnlxzkhHA8lRl0J6qFwaWHFaygVr3
EiiuLO1OJfcFPhtzgx7l/t52nzcVBKxKflA7jx5KY45FJuBivth7InP3INTu/r2QV+yx+5w37bhO
8eKIx8Odn6FmASfZq3p0Wo9HLw2MRboVVVqP87veqNwqMKk82P9yhDBVCZnWnDO2bK4gRkqjBEQs
6ws/IoAmwLJuXJGSAUgFjXFnmYMMfcqkuyndStsFEna/RiYAy6YVm8McOY1aPnA3yB/avJb0FV8U
Y+9onpb8swlh9CtxYd5dPMTlpvrjZYDzMjQgaj3CZTLHSeBJ/+gEhrvrV7z3JMdeuPgwyYwkzoeP
VHXWSomTc2YVANd2+UM4bspiyEijAq8mvBmjMMRXjln5+zD5SqLpWMBWs5T5AJ0z1Nt42z1/O9TM
rLpGN5EGlzL08lC6b8ThEKQ6uPL2fHfNuUAlXpmCg0n093f4EhnBfpuiqj3aigjZ/tYg6FWJ3WOZ
kLVF4iQR+Hf7J871gufiosQjKFXEWStR5yG84WtApDsFxDGAybUgXkmcPFRA7d7HFOPvlgZltAmL
dL1pLHnGqEXLvlsh7OWYpeFimZyVrDsZqwSriEED2jZ3lTIHWpwAFoNNmN+ZO26nbML0SINjOYuy
TPBAbWocJlgI7mkC/neP5zX72Ldg+1a8MTMAkG95nkP+RovxlDzRrrItj7eecVHJRD11ZuPEp34B
bqLJtthNx4ag9+gXH5w2MOO5+0zn0sxXM0uTebHbTsJbZzLBBHyjN3i7zhU/WdQ0jr1MVRY4bc22
eXLbjhNd4gSWJ61ddJbKV/qqqD1BDk/dm4FWIf5FZE4VXov/02+QdRdy6OiVnl5WHEPOMqfALOe6
dhn8PyzYZlL+iiE4ZmAd2zn/zdew0wfMwRMNEnDUOG2bKITZj2uPB3wz0LZcYlxscS6Y1x5jwicH
id7tmlTZ1gktVQyF7MlghzzK3uEJedhWIo19teQCeNXDzEdQpUtAfeBjXL/6cUaQm73Nn9banCFF
efSaexIjgK9VIxEtC+YzKJcXfecvELHcxbQrS5ovOz6fsvtBR3cwN/pwt+0qTYGf7mGT+xaLDeGO
s3KawtRoagR20HCBjJyQA3QCJlHpMrFa6uOyYkEG8iGYcc/FGVgKo709LGUjzkUUXv1pY4EViBdE
3kNdkc8RRc0UCCWnflhM+w8ZVvS9q9lrRbVA9sfZ5uK2LxtnUIi6MuKzmjGwZIWrJZ9nnJsrInuN
cQUG36D/EQZPBOXQxqnls9GS+2sPZUFlRDSD5Z6Dih89XQG7SQnJpaOzwHrvZ9OpRSU9vdtN3gtt
eC3oyY5esQCE0G5uKHisAIj5IiiGOL7AqYW0qNFZBIykTAUJUXYNEkqQgt6oT4Ma+dg0rW/NstnW
KXCK1N3MEbHW0WtdXoqwa3hDHlSWQiuuMnVUBDHepJ8vX9blbV7UdesHs5jUpfDnjXy+7z/+YAts
pYCpZTQpQ/1yLeKq2QHNc4BdzuFvJvfUYPUd5Hmk1ahWRTpl3N4oRIvSQ6pdLfa86L3NqTJjgHCL
rRkBz/GEbjwXQRd8rs9jt4CWHbLx7XC9FrujDSIJ7jibwdWeyW92eGFfh7dXjNgO2CNS8BY77C9n
mMOUGixZyrat7j5T7hZxzhJhs5MyzdvXVM2aDLiF/8j+lhckMK22uvQe2N0nG5ExtlrRwhvaKj8T
I+HLArnkG2oZalD1wjX3Gdp6b9T6vhSoB/OWsFZwwtjDbWHy3aV+RsCYWJ8xxHaj2e3vm4xv0VC0
SHZ0iADCE+MTgsgH2pp9A8AVyEHjqDxuUDAOuqqDO+HbaQh9ESMj58y6BWPvirAwBj5jrnK66OGK
UgA98tgRdBzpWrYwgH8BYuj3CkbIjPzkofePH+ChphWf1ary/zLMAGN6axSoid/PFqj3G+42BSuu
ZYxarJzAkf8xJHrVPLolDAzMdun3ip3+Jy6TXLTOZn0KaR58u5sX6UYzlovurXoqhTFeK2eRBQBX
uYiHBKiwr/qbY6ojSUkC1U4EoZl1xLNRDATvGomgLzoI44jgkaTxDVcSO++a8PzL3JuXujYglwFQ
3OuRldIpS0mlOJiZw4ir+2iyZzoJIm/rNetlzXTNN9UUAtUbL9hMyuk2iC4U93BqlIvHzxF2WF6/
t9GXmB4tw0VsS2apxKhAAVYFWnBPEQFFry4iKnGbGcrfdGL9k/puGA3SFN804ruyYJIvbZNAjVjz
nVywm9R0AdXi4yuaV2HYg0hQl+dB+CNd8gkFaKG4brRmtWvSwDz4IwZd/oPOtr1oby/lsWjSEv1F
TKA0VUAcy5o2NB1EzrPmh919UAlTqXWyrRcMJkSUEodwS5oVVJlfLrnbQXmqn37NephhdgHDxYej
VPRGtO1+BA3YzrtsKC9Aj436lE7C45OzWThCdL/5gDQIPeSFPSq5HCywblRZ32rQLJTGjtDHDYuV
B4RTSKdDMBdee97dee1fbmzydzCeol5Ym2pSVBhx+AvuJuuTba2rLIe8kfXwloGSvmEiArXUgYL7
CFDyFnxgiDFz1YInVYcTjZTFMs1urozCKo0DURIut61V3MUx9UMyTH5njw/sTCHmFHnyvrttdZpd
TGZZuEzE5rNI4Of+NuY53F/+7UUeTfwDvxMsMuKnmGSORM7Q5Z/FZO1lRB8HT0b6GhJhXh37Wpog
vFA6pj9CkAq9OG32x5AnHQOm4WURtQvKzUItvDSfqa7GLPCCrAc+FMbVhVc8BVMQQOMHzfFv7jIs
qm5KvzAKMGMixAp1httOvc2KWWjIoVuTfIt6rDN9nWTxkmYwMjrnWrR72CKGYQ/MDKjQafNOyLOc
V+evCOi5Bj0Fkc+iBBQlLmPiYCxy9iLT2Da1N/+b6OSTXNoTtZitDEwTANdOyaiEA6smWAS+x0xs
qJioAlgjzsuILGI0BjLA0U3QNB4vweN51ldXQkJrVjci79GF0qN8ba49wXUBWyvxiFuMVx7o4GbA
JHHePpDF8EnfG/rodNF1xCcIoXFwpUGciS4SZhiM6ARzn5ivFKveByBNHLjA+J8J46m6c1o0Teno
4EMbk6SuTfeSSuihUebUQh669hrqYETXwykFD7iy2pGX5b9Xc5qOnkZF4+YxyO7uAmodWsArG/DR
hiseTpJrWWWajDcRfg4zIrSqePau7DeiGoPjCqomutxxrkjVYE73FUhmigfWSMTaGo5EkD6d9RDr
xnqFfdQbGHzXUA9Z15A/7OiQ6Fkbx2d+HM++z7sq5JUgSCRPhhEa+5G7Tn85dp1MWqgzIWg6mO/2
17/ashhBEou4AelyZCJ1KQKzhzpeDhEDVsUTJzl51X5Mhc8HOAtK/wBzTv9sOwyENp6g9DCPoITT
KLI3ZoQdXwCohTLkGyvpurEB6Z704FnDkL47vKY22sejg2GKKWh8wvoA7Y3fOs3shS/bjjKp8UhP
BVZD+O/wI0Hv/iFM+LGy/Tjiy8KRjMA6sbS1uYINtnsqFkpiCs5XknTafFPwbknAdMXv6/8U3otv
9nU26thetaabwLBNwCqA1hPvYJHulaHsUeZ7zutzBlsCyEWHcpwetNVQ8wTekegBOfk8G7vifAvr
3fufzUmqxbH35Yyvx31oNix8LjWyqni5YkwzkjUo1gZbzt1OXntieyNQCVZVqFwNclO90vlz4cCe
hPlkHsepOG9CaW34r5Kp7ZqyceQoF1NGRTOHIEMFuX3H8tgk6VKFp8vjDsYFk0Y03g5YofdAvq6U
fhY8SVmjpNuWSsct2ASjNP7GOld67PPOVWTYrbNjn0NoYe2/FIsHJFWu2vA7D4pKW6Byxa5akAN7
D3V2vCBHui0cYS21whMEoNODQ2IdEyrt5z72s1hP3GrFDRuB6VkdsTjH9di++FapH5EuItV0Lo3B
hgN8xzc/WNX68AZ7iEVm6tfMIqZaqBle0+CerpcV/SbIXFrBbd6CtGfa0rGF6TBWOYml66I4BOp1
8AsKyZI3yRIsyZTFHM3+LCuOjxNv9ERBlxxvg2RFkMrHPWB7+fjVPACrYsy7ABLB+IO1Dqyig7XD
3hNkcjW/5Qk2ZANSVLCZY/9He4+1WHHRGEMPuvj6BPeQUVKXTJCrlLqZUhAT/J7M13TCGUMMbR5I
9DQ84hKplXO0HvpZ0naQkFflXfi4mX6KkNMpumv+a8kPBcY2aCI2oVHRcgbQwRwbj51KTUmllyRC
EVNT3oiWl2pTV2sq/HqYptpuHU2j/k+ACze/lh8zJJfQKq3//wEhkNxaUHr8ILzmDEPcBCh08NeK
8S3KUgiR7nih5JKdBx6XOaYWWf9RauBnKe+Q3lAhOTKux9QhHIU174Wi8bA9/4e4pwgaktaxNsat
ESgOEB4AfAP9Up1jExTgBy48ehi8CQanaZKxjrxA33O/Ii/SeTiYINMhZu1c5Dgl9A773qhqW2on
cGEs0KIKTypt+Ic9baOczUxHIkX89/yHkndsyzlGxlpOgbDMmmD4zcQfmCwF8aPrJKz2Jc28+dsL
dTatXJ7LFUUZIKV1cMTklyysV/RFw4ZRhGUli8nQ92EPdFMJj5Y47XUelsYFcUYme5kTGAqaHk47
auVtSZNpGrA/qx0pItFD6TRShD8hKLJFTFF2Yy1BtHK8Zuj75jRWbeze+WpT2kPwGqdjwTHw1cte
GaF1NtFt7AuwUtS7CbsQbO4IfbxBOwmJGE7J4jNieQQcz9h8taa/uoxC85JJoA7jU3q3BdAeHYCl
ZjK/1mUT9/8l+07kNtDlSKq2ekdKT8kgq00YyOtEMA/vAXt8SPixmwYSSMU7K2CjISb+fQByZAcw
T+sCQs4xWnC2+oAtHQ5GDEMij5646y7M7nJc0R462LzRMAGPLgU5Lqe9rmpkTQt9X8ot78h2yg7c
ljr6+U9X9ftAoalguMGvINr6FY8OKnoiljbo8iadEXBuRc44+proMbIG5fUXJemlMCAu+twMa9aM
cE2HLYaGvXg1cj/HsLE9lDWBd5peGfylQnlsr+iqTfe/fiu7aWwUnbKJbFSYN8j+qu8Se2gSkHRN
twGtkmwLEPcBwdtzlCKzBSJ3NscSEnwn3WVnjYSXAd39SP19x/hvOSjrQVtgGEq9Bhn4zUiDv1a4
SCN3DH15kvms3xZXE9E4w1tJxBT+IDMh+trDwJkhxqMk2JJS7Hx/ab+V8zcShrJeXSzLE8EQxanb
Wx+EvYKtGgM82OQflVdN48Y4e7JDAv4kiF1McSmf+oicpqzvPhP1Mz7NFOk+dmM6HstUIr7Gi/N/
Bv4aNvGSWkwC4Gr+PFGLGP9kBM6miNPOhwWP9OPZ/CIea3T46xyUhs2BJCr3Ws2fij2iYQpGrcu/
f3qZC47bnXjk4O0EUnFS86cZUY7dzEDw//IUrPe4180GDvmJXKX5/BPbO08nog5e7gUO03sTBohd
afZgIE/T3qhvXRrGFf34Do/nJu2OfI+DLHI18fRoyloMTSzC7Kz89fptd0OzGNF8xiZKz1AHOr3/
xESamM9Vy+b3OfJ0iYSUYDXJB3IidFS2A7bj6yHb49SG5E1dTQiXNYtIhihWH8jXFhEr4G8Ta9ul
tuSwcXOS9DImaDBfxgpPNcTzztdN9DxriqbZN0JaopZaURIp4bgGcixx8gfeAFU52yJzCezdH4vZ
1Qe0qBPPw7iSxPwNpRSNItWeOYUS5W94cAykU72o7FNQ4AQyRmMwkUy4kwTpim2t5M5ezZQXBBF8
byhr6cbUFTXeA3OHRzPyXndJsV7pML8rm8AptJwbfiRnh2P436xIQ75WldAbxgStqDgLgUzWpv8N
brTZ34qQbc14LwXE/+e4x4s7CGnh0vMj8nMczcASAAHZNFJ43tv6nb3Gx4pn6viE3LM6jIyin7mU
yOlm8Ibq6YpHq+bz3vOxfwUwBgMMGwbCd/1T0ngvynAe3Ed7rNXkfjInj4TEuFXytdxYZTPtoR8U
VGWGpV/F0/q+irsLph/J+nsYOYru+AmtnHwr+TnfISW4FYs9GO2CHlL/E0SBsvTmkTtqEjaHSE8Y
A6Z30b9KFAl4l8O1sffdSiyfBw2Y/ksF2rMpxWU93apgo2XlzzFTXwLBG+G1LG1B8ws9L9X2lfut
IZJss+Tie9ED7adq/KD2ibBqUp7pJwVOdOxuLX4J3uD/gpyZ1ulqtJpn+nUmRO2XebGo6UjWPsE0
/+KVVlmAdWBs2RBUPVELEpiP6ovSv9UI8SSPqfjMHyRItn9CXVdenipVjnt2vu1mX2LPc/WatU9i
fPwcxI8gCewWF4NEsPreL09eTaVXNy0QapIZF7Bl6KZAKenCX2gzUIQfErdSsKkT6sgftOHf3X2k
7eirGH0O8/Ao7KhQbuMADKvqriXL7F1Cbu8tm+pIYIBTB9SonZ3hBq2LV4rs+DPOePnSdNhGjK17
HYMV/gjD3x4qLN2fSOZo2nHfmg2jw6jTxqFSckLZWLCnSl3B8docn/rcAG244xRUR59Z18l0hcdt
Z1fUTJMVWWv/7Ji88yTEhiXQkaU8mrwCZLQxvuK4Xwpt5fFI2jAP1TZ+cJ/0EdpqSVYB+CfLUEst
nKSxaGSMINpcM75msa9SiCWVbIlmRYX0viccw9asJd7y0Q+5X1T5Dx7ISfwVCsyhMnMsjryofAv/
YiKdYHfaUcaM6r/vv9y3k1tSUn+cb83c2916YRCjLK6YFhXZ0EEOJYExisCy9Vvh6W8dt3hyE5rh
3NvstGJQXOxZnjw+4k2wG73cHWBBft2eZxVw6Oibmxcd7/t4HnCgnXiyYVqrrdDMaYodiy4LdyW8
M39sIm1UUq7eIF0dMRk2uvB2Jo6v5JD3Mtjh5x+qX2tJim28n2vNWYJH4xCJae+g4AcG+nE0NQNc
UhL5vtkisjAKI+KsJR3Cf1msUUduK351DmzYNUT+9zGuHvmc4k9Fm2MEs/ppAHAPEbmKXIAcIWbd
44qx89Ai+IBLMRL3Y+BzZX9TCThbjRncCbWjApyU+wlCUpUPCL36ckz67FrmLMS+TUpDN9cHgZrV
BiIzyHHjOKKHJFTg/MFuv6vCLOUm0MLBWeOGxtB8fnPifbf+qsBvqGoce+DFYHKcYvLOnz+JkXqQ
9kaEbWlyC2fYWjL9eJom7aReS2EXF5GWu02KV4+gyNDJLtUm5U/d533r0NNu8YJruSl3ZC7eg0+j
/+Q6D9DOztHk8S6JqvxVSP8++Q21XsYfmmgbckkJbNU7gXUTbZ0i/grLFysfjuJFIQIr2RykDc+c
TUUBcqgNXPx3dW4UgHQdlxa0vLQ5DbY3O+Av5EuqowisMVFgz6nzq1SyYhJb7tzgKQlVEgHuTYcG
OVl9N6lnu/q6nlEeDY9SKF2/dFl34C7N3/f8pP/08/t6vT30ZKs9LBsXefzl+txWP+k2ZdlZou7o
rNSpMgGwbrhfwhZgdGmUWPe4KUvPUld4ZrHFPo1vH/ocijLbLhajqm6MG5+xE+Xpes5O0nvQ8Ai1
SeNk1xh1YczmeKvUfGzN99+gHFtXvDc7eg238NG101/Kj0bbXLJp0j/s3M9LccjSpPOBkM53QOU6
aU3n7XNDf4RTrQMiuMwPe9/p2JVUCzzfDyme81u9qvVAqMewyKqjWyhD4h5vFNxhaAmq43jbwHIp
o68d4llcSJ1+rEp6pkyc3YlmgTPCf5A4dbWPl8lqWYFiOcnwrB6341ngzV1J2O7ehcQaViJn7s1d
WtX8GxVtePTZCyjfkSNP50mneC6qbESJHliaBbZjNjvtPN27Fp/drnCd0EdZKx+UfEr7bHTSEtsk
qVlV83/qRgR5/052uP6fnWkzglyAZ3KORuN+jPrd1bKLlFgMXJQSSKCLBIZKdrG33TqQnvDgzIUg
GhF6OVqdxPN6Rxusd4KqB5NactT4i23bswjOq2wP1mrGvjIJ/o7zVMoZLAnemne9IJrwJo5VjoPJ
F+PHBGHh0yDZGt3v3yR2SrHvkdcysc/oYbJLGLKF9daCJgl/j6rmQi0Ad6qMoC+Z8mqTHkAosM+5
In7FQhnwQGC1LIrlMXn7hauZuc3OcpYju5f1rhSn1L7AUV30d3eUS5dHv4EkpGxf9YAqiCH0Czv+
XtzkZ/JC9sVtiXVEoIB4KUZtYHUGttt8EI/vwYhI+DchcfWfvIrGV1gslWnjBlAaYS727d7ek2oO
Znsda54s28cCIDZzu817j6RdukFLMT6/BFEFdDI3rDhd6l9O4Cqjt/eFbElTq69pG7hR3+QFmwDM
EIgdlRZOV4t/hx9eUBL5VIwL/59a3llvEyQnIRjIET8N86vCmjvlc7HboqCmZRRMiBgM4yLSPQqA
xoMaWtodk+HqB1y4Mf/OoiyPkUyF74XgI3fp/PIBkPzcDDo+0W46MvYGOOyKy04xIJVw0QAvG9eq
CdzYsyqANY7gqM5TaQ5USOYw+DhjP2WpjcXbpqMh/u0/Z8liCJhBi8ZMcm3KoWbrGzuvQR5vV0m8
dbRoJRgXZAusr+/kPzphLUU0lXtOD+WfFdDuag1S2r33bTOloHSDjzHfnsUP6Mrd346YJk6I8Xvq
egqa6xVSDvATZheF4PxqjhC3946wsZubqiGxg+u3Rl+KeFDmmnfGq9Gdmk1orhcsijP1Mn/FaokZ
P7yyn2ZIoKFeeeZlVG04qmf46iDMYMAaoxP2dazePNGD+H2HoZ4wGc4YA2KO5Z8pNvZ7/2XUMqNp
Rutfb1/hNVjj6XOVEqePUNZdu1zbDssM5+qK4xY2rZj69u+fNe6w0bZSno0xCWroWjDJ9e1EIpKY
7rE1L+DOx1MVP9KxfHh2WrBGBG+2BJdeIn27FnIT0zauv0IZxgaqrrYA8o77pPwZ6gT195lG5ioP
M/NYM4o9AxzSob+nTP69C/IgXYf+ZPMaHTlYzBh3WURViu9Lz86SpemJwNSmEPATFLcG5jH5EATI
U8LUy4nkRXxY4glrjYqR6f424OFB3VO1tKRZCXyrjzHrdC1TCH4SBXOVl45wi1+DpF8DNtxW3qeG
u++OzTl6ICSAsPbdnuPRMcE3gvrzSz77N6/KaXZlISdSDRNrhvkoWLIFuIcM312jYzAxBxfyImP1
2+UajYZpGmvxIX93Ox+IfSMOORMWqcyuZHfcIuo6OIjusXlWwKm0v8QsvV8G1FJ05NnpyoNTeM/V
0vCt3DpJQZ0croC/LWpcXYHppNTFt+RIWx5WIZDbn46NX0fspEIYgByZMhtaTpjYjL/yCoYunlT9
xRIOvTMsz0x/lg4gXSJA5PJnTP/0IjL2ra0etu/KMK9R384L/SOSvF4NqXp1DebyR35DUSRUu2NS
g7NQpluqbqE63vJRuTRmfKrmKeuJtF3uU9drdlKCxbG+JMA7wJIdJbdaYNJ+sO5NeaiWZbQeNjhq
AWlZ2oPNvxZyfYakpQ9F2JZIHljgkljxUYckYQh6Nalj9lVWErp/O6sU8zzngCO+SnjOYIlbMO0r
bfZXL0mLNTOx8eMEZCxKBuSwuTrGcUgwFEjcTB7Pd0JQEoXOoofgFR8Kj4low7xm1/lMK4jvgjEg
O8eQ0R9l+xyHa1zz3zMrLX2DUT1OEwIuZFdlC3KaP4yO/o5mNn9PqGkQsD0vtHypRU/NPfio6bnT
lY6wfKlQA7dc5AQM5zLyUZnoA60UHnZB44gmCMi/Sc+SUsPhgogsKUhtbr9/shdSB36BpiR9OCNp
WGoYvetKvaUEUOtVNKIC1iCvpdkCxAaGZj+14KNEQ+P6Lal2NN6gxJENl0bPLJ8DvH4LfjsPnWeD
UWaJJhYjRA+dbsMAO0WxG3Vz0Xlg5ZUOrupsF5XpF/ihSHA73fjdBQW9uhqnAkXrxXwweW/65xSq
mEdYII+FwrpwR/pd5IwlUw+ISRxtWnFEu1I/PlaxJAXJgybk4T+L/xLNWzrkfWO2UamlsrkgPrGG
xaoltnVjnsPVyLk+FzJw4A+kpfe/Dtum5GxxU3ZH/fObSAZz3rGyeO9PObrK7IbROadOUxHhKmO7
M4j8xS0hO+JZpDO2LGl0ZUeZbcNdRIH+VEiQj5ZWx4Bwx35MzWYOnY+v2hL5WNGUQ2gvBlqY4SdH
mMNdBF8uKNajZ54tyh4IF4mvnNlA9YqXAUoC94bMR2S0nH7XcpMEUs8SywFjrCZyVIjBTwbN+vgb
oISubSQ4966BWpkCeYPCq0FcgXs6pVl7M56u7FNJcSp1tSfHKew+3MbcejSFoWc2QuTzZyDBql2p
nL2AYeKGKKzjFgiiUJA3Bh+T5B891mdLLdnWXc2GgSusmA9H8gCuziCSKYh2fUkbaD7kWKlTybBL
vgzHL6EwYtEFFr0YDjWqAa8c8saw7ExUvwjV0RvMlQaqV7CQsbxJtoLA7imGHIQijgMobWFC2VRd
bhCs4+vx/4gaMuEJXrZmR868XG+L6VMrRH4w9820/gkyJ7S6Hg1Oh+tR6GSuw9/6jG2Nmm3LONzZ
kAmZ3rmH0hzTM3HD6AXD+/2/yMdj4PlAvhPFb5Qz5gooPWJre2rHQqpXRwApal3luBPvNDneEsFH
Bxgv+zI74ckktWHGepFSaaHXUBzJ1z/1EvmHj5l1xGT7lG2seinrDPcjvet+jzRxrNedELcpyAgi
S6/Q/yTiAGDSbJ538DXIjnKByXPzATJnsTWr8CFWTOHu94R7waQJvAmJwb8l7rPDU9GfVrqzYJOo
AGi88RLPqQf+ZV59hpP4PCu/GVwN3vw95aXLo18qFfgM5/mHpI7GX5And0JZa/LHLhtlvcadYK3c
88EQaArQVarRMGxbDxhvqZBd+5FGaOJE8nQsWU3ujNc/Bs2CqCD6kEOaXsmmdE0foIidB1bx26BN
DgkYr19lV+ve2rSoMIuPA0Gje9U8p8T44ip35rc5/TolvUjohCSlgDg8FUG1pYA3Ym4YZNX2KWLD
3j60K+q2DWtr8vjuqoOPnbyY1wUUKr84PGWgVmgvQclAqGe2zLnQGyGH1JyajhHrBC+VhUfbBS8W
wxt8p8wwsB6E2ziLTSmsMIPRNIyitxYsp3NnZv1C67I0j9KbPJUtQdW0fvHr8sZrASh7HZ0uqY1w
g4RgTpNZNwjLnTSiBH8ZJlbTK0br0exxzMf9iFMjBtj8YLqYtO4Hhx0S+0Baq2u9+lpHROhrb0Yg
ECZotF7MyoVLOQZNPJ8l2MiDnAXYDym23OiUxiDtRnlPZqB8AIw2nIcyQ+pUdLC/2B881xETtnFl
PjaxuSTFVMZSSpbn0si50Pzz282qluI5uWVBgTVBIPhzM6XIJJHuYX7zsNCQYd5P/4ixZNR32/KS
ntKMBWyzbwJWmFCrUgpKW3UbIRI1QUNbNh+qnneORikdcpyEFRa+VN29pFFvTqH6aCZLiPRo3pRr
LVP9eN3dVz+eW2gd+Kh7xVgjsSIuY9DsvmxA92N2mDPVlHB/JO8YQwZXdfeeACo9LGSpzDTTZnL+
AGb0cTyPg3QaSt5bZdv035xf6PuTaL6H/FUnKANBCaJAc4Iy1/CWqYwddXtE47MzFQ7apKA1c2uw
AnNOKZcmDYRPknsOOvw958gVKzb0k6IZbdBzltOJBxkkUIBt/JSU6zSFV0q2/kXZOyCXlRFi5sr8
LunMNLWgmjYoSojREIX+kpStkgoPxFBA6Vt4hfRcwuXs9UOP63kHzAyl5OmyA5PcZgtJ7pMo9HJB
DzzMJOePqVd1i/L4QMyQ0C/bLlDGnEyuapy27YiDDCOzn/UXO/p/1yMDX9K0mPAFJora7xnRy4LS
aZ+SVMLTkaE7IvVtz0ulzxztyWvIBx0oCS+Eie+VSlp0gKjfzn0a1g9CCDqUiHV8J6dBNRwPApi5
lHQeNr4k/MGcF0K6RgvmlukXcKdKltn7Dvvs0O6hOSslbZOtz5u7J6Da0ToYA3bWVUlfE/G95OYm
snV3Z2sMEys+qnZM2CiReDcvRgihXj10w+a3XfZRzmzB1Ysmkzbi8nPi/g3XExqJetqh///uXFz7
6FVAQBT2jrhJfX3lEMgC8kPjwfY8Ek2Acr4Fa7Ki7FJNu797ubnAJ8TQaP5UqDJNJ5WBMJFWpIfG
qnMmGB81bibB/Pi/SvrOi+bw+qPR96AF7XZ8HERcKRfi3dCV6Pn6mtgoMIZjTxaslEQ1vt5h2URI
Z3KDWxInNeB+FSlsou60A7wKBc7wegIqoJ+PC2kiKKJiDTihddFQdbiD8wyLNLGw67Bj0a1Mikd3
jepqSCIpVO8v0jUwS7nJk02cEHa06xa3Xo+p/7l+ROWiNZZzpnkRgA8VxmvTZyeVEcBsfSjmPft0
5NUug+vvbbzzA+e02aCW2f8OYz2J000uuV4z8fXeohievSKnPqvbY7+JuZjx2hxt+np1AwHqB7Ps
x7/ErxpNG6dWu+fxLsFGPwcNqvROmakStNiiv1BjlEbB95GyHMkqp58QKfnc1DR2qTsdc4GIQYpW
LF3vAm1u2izjO/gtyIt0heck4X/QYGTg5zOUQCbi4a3f3M7rC2MpZF1Og/liJAxQJmRA70laVbUL
qT/G4bdDCKHcL/zaRTKK4FWSw+nhrmuL3iZOKxxg+av+8V2YhgVjwltHegOPSZQOCW0wqVROlFlc
erEPNeWbbA64DUJgaTeDSzFLI1zu7UIriJg0jgf22GalpuUiF0d38GodGMv4DGFFgH48FnQeSKJ9
b+Zfl4RvA8gX65sFYnQpSYwVggWvv/hlbbf0OiSnK2f5ewDd+GS64ZmTMWQj9eMVvyAxlqQ2Ye9Q
/5ph3fAQIzTKGVVqnjCty1h69gNjx2GHUejvH2bpXUOk39NLVi+dz28w1mI0flwL+Nb78oDUL8js
sy/5fVt6H89LgAed5C/tbgHAVI0d6+OYvMGSc/L7WYIFT22eUamFJZHLo1+UxiEP5moJ3h+UaSst
Iw4d1FTYNfD8e797yD1BqeglYKyz6NtXd+yC4PscsHs+ETG42Osk+EfhJ6agVXX1OrWi2TrXv2Ec
rAxSNjj7lNZn7x4ZeZM11Cm5JkHkhWtynYpgB7+pkh29wZdgugD3psx2Oj45/frdpF9QmBqrIumy
5qApAeGE601oIjbQdwJdT+eQwPg2otvg+tLb31N7X929hadvQP2I0nby4XeCg1ldqBm8Doj47Vk/
hFsMqJVRiPXCI+Z18wHuEC3M3Jngm/1RifCrUJvs/wl4VUxRFitYQ03p/wYbQKzBrj1llLsRhzso
v1ma1XCSGN8CaE3fN/ux+0rjvrkbb4So32dZuBmDO6q3HugKbWdfLueyUMs+W4QQyky13o/SpTfa
Y/+SrO5QEZlgxRXEZMgN0n0xrGfKzJiEWGPJV9ghE9CX4GEgJ6O+h6+4lrVEHtWrJugi7GDRxkjk
AGZQ6/GxN6xtNdnsIa3sOReyfvpykNCBOeGYYZleW496PdEgwsE89k+uSviExTDOll6DMsi93GHt
p/o1SR6ENUy12rNdtPUV0ciIz9rTq8nVYYW0qkSNdlqCLnSwe3kw3PzVz+o/wm0H3F1ttIN/TT17
jYuDWw7m92/XFoyXxmtILTesWDutUcd9vY3Fj1OgRhDQUkBmzgbHbSCwVle/vfq66IPoj8oig8ZN
uzn7lQkt6kDB9j162lGI4or8ZMvmshAoAb2/jqvMt1a5ye4BNDrG5np52sqPCiH0yFIeX2aJnsIj
X/R44BJzajtyguYF0z9fjSDL5BE6lbmY1+v4B0O2NFQDKMqrFORTeZ7iaRf/8bC7mJrfZ8Q8H2X2
pKCZJGxukHjiKI7hR0VBrafwnW3wXD7DiKdZuvdCmBUIOoWVzGeyFgJRoGXvy3Wajci1wliTvPCv
zClxLSo6p5UAtGMTP/+KVaynnbWH8n22IkDHTIO6e5iwwdSconlSfWqrgUaNG99WNfSSwwNHCjDc
y+KzD2MEqss/g/CEJXqGyPgMd+kDG9+xIqBr8jdCzHM9rFHRgT3XsSu413daGrKBJ0sa/WmnVLiz
vJqu/W/1zHbqWncxqoMTvX+GMRzt8UsOQJsVy14LkrK4sSpKf9v77PIrxtd0TDWzpqpO95Cr3WG5
VHPQCav80f2VF3egEj1K4AQ0rphHurhv08MVXuGYUGk35xg34ZybA5QmIIFRHSpSqodnIMjhbwTq
xnvpRc8mL7yTDwlV01wRE2INMXrR4AP/16+uLnpFbaGKcRRsoNQcDLchQzrH12KwFYdIt2blPLCO
aQU2K/2DFM+HW4ZVubui+lnFK/RND9ED8UdK3KoelEeuKCIpWF0gwGlm9FHprdEQBM/2GgZGPYjC
/LTz7Rgg0tiKxcwFCTKAmgOAZQHjKfMAfrUxyhx/giMhkEPpb1dtq+DoZEjI3vM2qDEu5fWOfrjQ
TUMVt386G7Xbd3wz/2lCpsJhEWUCrZsu4k4sItC6WgxsMAkgfJ3Dr1NX67m9VJOOkdH/F8vE8Pvm
+TRza9ah4iam2B+TV5aZf/+siA6qP2tknCXHkL9FxAcSBlIPKMfRzGgGmDgRRlNKff0bnnuKwYSz
eS3PE/n+woiRcgkiQpj2+sMeSl3xtEcqwRlcgHulCtAzphPSm2CEwdol+xtC4EVsnyjxSkz6/Twl
hfpdlDfQWUJbRcVavMoYFgErvzL7b3zxb4DmQlVF4XlZb2BH8jaTximTcjwxQGE6yA8iOnyaUbdN
MG7yHEKk+G0l68EMSTkWiKlTvenBM9vnrGm+GAZNW8qtJ5egS74pbJ16GfmKtBTvehk+FA7ozwt+
crm7HY+CqtZPlWFIErPRwwsa+u5C5H1uAhnNVIYK1SOSmz9S/r7UH9n/pXHsv4grigubV6HUv/0y
1975f0vFFvi8euE2yxAAwNYMNzLwS6F9nxP6d4FfuujWP+mSY5xYlWFVbd6eMm/PrgLrI6b9MxfR
G7kHDg1nCJUofxa8RIUcaOHQZ6SMBnZP9uoAsrnf9rLL/T7mrgwAR1QSgtavcH6M6YUDWhvkDhCn
2WVIHU0aE5Tgbz+UtaznFLxXFcNfnYFO3XChDLEEHrWK/IrBsuWI72gHRYE0K5Wd9D2MLHIS3s0H
pwDFdUxaFxVUZ1xtBJCApjLlF95DuWsnldt9OKQH9s41bEsPUY8vSHd+jMKoFVJalKFsl34fCo58
pqx8WiPyFiNpiHAfTK5ulk2tVAqfcYYu23Z5Oy6C5am7j6crt2kW14UfNZpq4oldnfN0sqU/iqKl
GK7rutlEVfEKPG7u+WZHbxCmwjsN9IWTcOsFt95eC5FM06xxU7kFHtU6VEEJ8/4uUu9QMerOoSbK
c7V9NSmcVHG2YVJ6sRIwOmGogtWhc70COgeqD15XLtWM1T0Sy2uTKno2gNwBeZZgdGo/Em1EAqMO
bDY5AbXJD3sqNRzzrFFeALHr0S//WgSzeDYenVr6Ua/Qj4eVW24NnijNLPtNXiRS/JxTWMRR61lE
9ZJu/F8e3adTUum9StAJx4DhqXeiSUlCk9nMPB2VSqldFbP/ehef/7GUEk0rdixpu37GRD8Y+69B
jYJBYrUKYrn/gm9tGYGQHg/IAjQawjj09LClKJ54EBtJy8zFEAfmKXtBd9AOrdvCxkGXWJ7kuRa7
utMpOacVYwj8ioBmVDkNhrM2UXLABbymCrGV0OPosm0Tp+qFSmfMBSOcDJM+6eW3nxJP0N0QCKBi
EV8H6ZeDADM5+V84Yeds3vq6U7BmO/GmoRa7Exp0wdooVu3fKgIsMgdlIKP3BUFBQLXaDiQWkJxG
VVMyoJdMjooMrWO156FGII/n+qScwz/SLgpQqe0CIoMnEwrxKZ/8Jheal10o+Bp38MiTZWLRr4X8
ELQHwQNrZtM8qo4vRgjIuMT5ne0ikZ5xJP3vEqFvU2vl7zXL9fPUJ2MZ1dCzkNl0VfCTTn8HCSxu
4BtXxLTl/1K+gm5XyP2n1AZyn58x5RTJYjG2zBK7rWyuTuRKmZLjUg9rbiJg28PmY6BPrCBvzCQ9
Z9p6r+40L19803h0kLu1VCAn8uqg+1gq4g5yUu6KxbotOAXO3QQa6S4B3KIp4Ob7LHCcmpvEicDd
eB4gB4ESPubEqWTpK3hLMtmKAEygkD/9Ot37+wg3V5SMXN6+rO+QQoRYnL8/NW4MuKrhEK7KOBje
Q3aEA9YEIbKCYvxpBW1mwKPE5zi8WYZhN2J4v3Qu6sTH4xkWmFOo+i9DCjY6QDXMLVMuQ/tf6lLS
evrBY9anVM1YB61Zcqtq7j1fCw3u6XFULn09a0cT97RJb2QyMRXjER3y3p5JidYETgHDj3OBHuuB
5vtjYs4kkMILXqzGsDMDoKsaJeWP4ihXRuz0I2F1LzUW0+FbmvYuvOOhBi8GeTfUPeJyxSJz4uNE
dC8ufq8Of8s3Dm6HgsFUn+Ff6SiXi53kDN/MyXejX58I5azqM05sg2H3oqhIdVw44SrVTXMRSEkC
Nvg/ZCK36qzVTXsZbeAApJnzXjVvDF6Wbzc2k+rsJ0ZiXQJC/7zfLcgI1QGsKYwWK48b+Yzx7kHZ
ccfwe72orsANg8rfec6mhjuUbTCy8Z3sqn52DKmA5tZwYLJP953QijPz2dzLcFRO28HLkxdFarxq
KUUqUBuazw/yeLhod8qxu+LuXtyaaj+uDo3ugtQrMtwmr7IZDqsy63mBf6/1tNi47WYK8zOz8Dnn
hTzOqCtY+Wl6M5CfafUNpMSmDNAoj3t1Rm/C8NdqZeoD/5UM5ZGLSRtaqC8PtPvGP8l2PxinUGTk
EDJJQBEJTvlqbMANLqhqpt1uDUzS2DG9FCFuy/Xb+AZWcE2Ja1RAW9FkEkTiOwImJSaa9PUcDaWA
H5kYKiwOGYczh6ZsIp8CVjeP+Zh9l9UPC+vyZt0edlMi6Xq0DHGWd6xJW3HRfAJwQDiW1GD2EMNz
OoKJGLhuQlAjOoX7DG2vr3ZyJLZW45Cg79w2vtxTFPHnUIQBBBZQycPrmZcWoWIM7wBpUI5Pzt1Y
xPOXHU6W1elQUCNoMygyatLV11A/Ty1sTjMe7BC9wtk8/8EJTQpnnGHy0gAZYrHmEuJM7dQ3/N+f
os/0qblmFVd3ZTqnZxM1w/KlYl9bUdgSkaDAeSl/0iUd4ydu8OGVSucwdhTxDOUoIULwycTLPVQu
rOnl8oqczzuk9NxoB5py41ftfwFRSi5cOpNv+PKMAmdk62GetPQ+dxEKs1nxG4INOmo2ERYfntct
ZdFKoPbROkWdk8hDjhjvJFz7g3DPc3DkU9Q40gLF81n1X3CvglBWDJ3MekAgZLyarrCtVypTi6VQ
bLBb83+xemgUBX21sXTa9QvkksmOQf1oaLys6eJbXVkyXVQD/1YzOfx0wa9/aumQ3ugepVqMwaxS
7AD1XHKDvWofZPovaPlpYJx7oYF9z7kGpGSUiUeIEI8V5nEd+LS8wXioczqwUf+Z/4+fKjoTfAbN
QA+cTSZLDQtDM+jGN4lrNKEc6KX40KrD2SvS+eR6JW0EjO8nTEgSpa+YuqnVo6oMAwPP7pzZ936v
Uf+xmtG0uGZMlnEbeG0Vi4en3mguNx8ffsA+Vt6/bPBT+ZfAtzxz5ipP532Q2VRgr8KDnp6UseMM
aLNcWn2Tr9EsNkpvhJJwrMh9R0Fmoflz5LKNWBVjC+paevm5L92k+vR2jRsIxuQXFxC/dFdgxNKL
ZMn0wPE1d9VQeHzatgJAXKd0WiMXS08H8uh0Pn9Hz4oU+f8h/Wo/f5UBx+A/C6odgm0j6Hee8bNi
v/NmhxYH+gbMxbT2RSFoBHVZQQJlXEOuXnVDabeb0iGfN9TyHr5m5ss3m5yFmXLj9GQMaz46byNt
4CYPRFoAZzks91mNQwh4t9PwZWSFCFGfAn26ugA12GMnD33D4UIU7OcMG0DVkKrrB4x/+C8sb3/i
PkJySnmBDeH29PTazFJoEjhd+CRX3ljKYkrbgAoBfJC2/zNq7XEoiA7oQPFCQBup/ZCKeoTwYa0v
oi0+q+sA3/cqT97Ka7a+7SFHYbzkxw8NMKruqSTiREIXB0D7MMOzAl0QPpPyEMvzJWYyI9QZGSSC
WGDjr9K2RLuUH8OstYskHlB70U7QkA6M+Fc6f12SqKShWTD1hyqyWI6q5oUhDPmVHGfPwZ28aE2L
WBTdk0w0Gq+bwskdJw5QzGjyqU9rml8O5upL35ogw8ydtSgNYQ9SGelpeC4On1qB/vE4BWc5nwFt
z8uC4f66H96LY2rzD5qEpdeP3wiO5DDBzkcedYayfcKZYuSaseqomgHeDf77tODct1uSpdTodbQ2
t6chPVNCntBKkI0MQzRcrkqZFV9K7WPSysNtOtDNoYT8qjPlYSsRemxIZGk/N9F8o90SN1N0cR6A
gUChSFFeQGiVHtBqiqiZvIfQ/KyWq+FHfuX0W0IO7MyMqF8Pnft/4uwC/dMFI1+pOaP5OjB1rASO
K0FySeB7gITndME+2I6zIYV23a/Y9IF/clpMkmzaDJPHdQeU7EyQhrPmTD5QjS4UkgFrxcwghobB
jfAFJxytuqoh0qeUKSZPyCYKB2wStJqbjOqatxDYGRSevPEV2z776JSvNOqmBNTmYxyE6HK299tV
HepJ6ChyhQ2F0H9cGziW3ESf75jPFAecANsKEn2/TP3GPQ+xMxWZfRYzFsUeeQYMUVG9CZSXpxT5
ukVinektIwen4dVX2ZCNTNefZWtsHI18OgumtBcZ96P7w54QZDf8YH+iV8DavIkhhefNftzoIWn3
c0eghv1Hr+oPioRyx0Os63anBXXDpmFDZRTrq5FhBiBWHEMoxzrppc2bDS85Z7UChnqcD277peCy
FBqsApaWrHJqsaHRgOYR4O+DoCniQwniY+hpiUnCW8h33FyzT2iVCRBrHMt1KksjBnvsYZzL9wx1
b1WewbcUPLnfNH5HrQad0AfM7HLPXW9JYJ2xsp79bikgByfAzKdMYkDDw4EyYz5fnNMKFMzHiny6
ereIiCqjUSuXREEeHgJh5ORRzTh8XbTiH0J92Y45MydnHbk756Js0xGoDa2vFpefwm1okRFO2Qxd
2FkKnRXRoLHBSq8lTyDpqPMV2cEQdLUU+83W6o+im59/VfLmFwUXFvBVYUepUCOsOlrzAZgblj7s
huARuIMLPiJzlneMMotOzKPuWg+fYFZEE+P+dhMryn4hx2wd6kazUxcHfRX+1FYilwHBzhHf3NOB
8B+vr1854nHYkYlxvFlYe0O+xcmnixs42sUkv0IS9y4KEe3KulKYNZG2AYy6egp8xvFHHgc0fikm
rsC0Md2E9Ble3u3/yXK1iRwicsewkIRpr/GLDX9sJVRiD5xg2otyE0nqas2/JP44XVqxZ0OGgycB
ij5phLvulMKVWPY5Zal8xDqb78qR371YoQohl7/Mgs8Pw1Ewzbjy8xt0z0UIVxKTGD0AIeReS/Uq
yTy3+wAtXIHi8BVcVAnV/d5EDcXhtOf8+395KzdVPlehi12wukOI2l8IOfpj2tWst4ZHjXz6UclM
Oafa7hGGAqx+Mwt8kfEXdDcbDiuTGZd7RI7C1+vqCVmoCpsXFPf+lAhQLSej42Zw8haiCu9b861t
C8JNWkHWaWRpXelwywgo5mV0++SAZWyzvfwbfYjP4dl/U2NiLY2vyWrCyL2vke11nbVMZ5ew/Cho
xsbcHxJOsBy10umvq9OK9RM2qnJbQ2O/ePPXA0ZX/aZtAF1Y0gl31tV0JEXFRRJ7VRG4ioDvGcgU
6TzUi8lwwJl9E2UWjt7WrnoSFFhMYumu2pRtoscsCK+D/oOaEOMbLbseWPIYU4mu6C3bcWUf8ZV9
Zpa8C75pILLCIpgjCGcwF0AJkZ2NoMS4NaaMMd1hyX7bMl1OLv7sPx7TayN+bUqe9goSZqZ0ELB2
nCQ3WS1tinARuFiPbwsQQsr5w6TjvkSzdNQXDWiGRWbcYE3vrwcLZyY80UZ0N5kDkdWAnZg9E5F1
kOoH82/dZXVNtwf4H2UZlkqx4wCc1NJJHuCJp5TeqTFkoEqaPEXcmjlkBEYXhsPqZzHV3f2HQHnS
Sz8nKiWqoRyHLlyiNjnXh9hWrgmzoUX+lW7FZs5g6OiLUKKgP86jQk3bZBOlGec1pxarP+Fpt5LK
7iNdrZx3nvFJq9nEXGGuaz/+KjpDAePHL7nw6G/qKCcXbrw+pCPvKIUUxIGgHNWdf3e/RiC5i9Na
L9eKbcf1SxyPEakNlB1VqdCdx6s6DkF3k1+Yq0E76EDZc7c1oqj4jfhNmlilMD9GD7sT2w8OpeQr
kTAEVQHzlCpZ7EXV5MLEuHB11UFIYboxQwSyG/qRFZpemTFOl4mDbLCd5fKLMlujymWaWdFbeVuF
jQJ7lD1vCiN+HNJpH4TONIsZzwjJl4h+DzPL7KzAPIiKMYe6UsHQ+6G55PRBIN+s0lB2cGvvPJF1
e/IJG6m5JSrUgUqgfauKF0Grq1Yj4x8NUscLvBZO5tMkk6CUntVfpFXz9Ah7C2D+eqE9KRj7jNDk
g1IF429KFl8Ql0zIdSyKsEyo+pmZ1SYWAE9SZbFPz8eQOE5chi/Tnmvo25rDYoHHqZjelTCdyj/o
1prfc8iImMr9slAjOjPdmUvHKAYBj/Lz3Wog4qzPLgIV8FUng1Rr/x/hGvTQOSKl+teZu31HiwKX
7j7roRqoP0epN/I3F6P6/IA7/rt2g6fyfBMeyMSbLXeoga5zyZWAccmfTlUGAptWBnFl5DUuJxcv
sijImib9ds65izvYXd0KhV4qWkV23GhCrBe/sVbabLv02TZaJT8cSNyqw08Wfc2EuYdeDqimeJ7A
9utkDD+nDkFlTXNxRZHN9B1lmG85aPYzKYx1D/9lC20g+wJRA6GPTIhYFGlAuMR8hTkaUsywwdA5
KusmqMSlzukz5tkjpvBrDc4AcmPwsK8znfAMtmbLGy/RPZIa43kI00JqJNUNhSNLEX5dRHEPbKox
wSkbxvpUngsov6x+8qc7IKKELhDzvamZYyZ1Z9HjCUAX+2RSPp7D6W2ol3ti1zn8RW6KEBxxyQ2M
q+jfUSsnUaJLnc5mhNKETDvXzt+NNI4kxJQBlzo7V0S6j/XWJ9JIscAhKj2WMREDrNelzyFO0n7c
qPp3H8InDAs/L0bxTSIUFlgo6LwKt3sMZoKdh0R14S86K5FjZ8mYE83qIq1qslR4oIHJhdfHyaFe
ILy7/fqtrmsPEx0zOVxrz+yx0Qu5/GXJR3hU4YUYnPbVv9EVDa4Iwip7IasMNyyxCnZVTz167qNZ
5pWMMteojZbO5Lwg14oY8yHew8dJOx87+NDa6CL/cGg9+gXfo4+wxDxA3QLdvZqtAmWTf2l0wjiS
3lcNVYLYvOWiAIL5vR/pOuLqWntb8W624VClY5HU+DyTGm8zCsm7jt3fytCHfr76sfokA2snOVaZ
nWFs+2XcFsKYhUuVjl3GAVK+RSduM/dF09GuLIBJ5Kuti7P05GY0ea4dKLDElOzWdocZJ+UgIlKn
/6ngNSqVKP/px3a9Kvc8V2k+ic/BnSxoILr9z0MhtuCy7FslYwBrLzTsvyarQCB9uHkmO7qa/B9a
8se9goIKYDrcMLbzR6xaza+GNUCNttH27j1TtT5glC0xAaTVseuKfGWprRHQjxZK7zs6OY8X3m18
pMLexjeWr86IkU9WrSu3z5ba1QUeXtWA06IghN1fLVOURL677UiOoE7oN31S9q+vVeksCzpZhVwQ
mWPCDO2UsUPwf9nh+44+mgV1hiiZTYWysK8WSzOx36As22YyNOGEHTHLOx7tiDZnZgQ1A8a1bH/z
tupiZcJk1392LqBvWyiiKKI+dQAzcRYP60XoqIC3GXbH4hDGom5Ppfxe+XYp4paVPlwKvUnDt9yI
u96BauDbqSFKzCkVpOoxTWVYPkWcHlXLFKscPo2t5PnJw7t38pw6jJu9cJf961poAoNo//Dz/1QD
kY7E2IjwIKVqukkxCfrT/gWiV1U2cDoBZhPJZAsC9m5XJidNxpnwKJVwO54p62OC98wDWOUuXNuE
eWVHDUhuTzXn6M9ZrXRKP3mXOJW0Bq+YkxmfEVDCUkgtUjNzKIbQkFvAL/QUcgJnWm0nYBN52Tk9
lIP3O+xqJR25avAZY1Cp4U18NdOPXsKo7HMB4ZViXgF++rodxlHiCeLuAVQ4SwwPi5t/Qc228bVR
63LoXVGy2sfd/enG8ePlrkb466m2VMbK+QjdKbagaWDbJi7vEvuLMXfzsTeovP4vL8P7kW6s2jJf
EcHoX6doCf7fUadcf7ErTOGfe3wxbseH0o3WaAHF1tnNBPksFfkFh2nw17CKIvNIQLzhslE74ADG
gLAQQRg7FG55V1XMyVcN7RWjgWWTWgyzhHsQvkz5qDlREobXVSi+xTvnffDEObEclb+Gx5mFiRj5
TyjprO+7K9OVmoCh8D+zF2A6sv9sKCZ6ZS5Ko7sAXJhA6oOB2wnR7BGhNVvVx4m9QEyiQXbIlo1O
guZ1Di360fGghkj/KtYg3n4yzY/pBoZxYaYJLRHed5G9B081Gvj9Dq30Tu+DwsaxHV+lsK4hxc9+
KhUdTA5Ew/FpofBUzibpS+XAW4Yo/87YF0zStsHhk1nhyYvrTs0cjEsleVQh3uPm9ebGMP2LagIW
uoKNH48aTyLxVme6dHpiFmw2tG3evuocXha5IxMMh6qkjKdYsgu4QSDOFanyHMcS/OgAoqhPj6/f
emdg3SUwoxGuDCuGy5hZQzft05LhvJXEAQ1UU2OpvW6TZ5FtxrIMha3FPaapp1uhqMK1OPTgu/5e
OH8p4H8gCirEa96oYPXJeaKETI/BSMEf/mfjDRVBRgO5o1XMFhJzRMrPpEZx3WoiqHuJZ9hLA9gx
hg9MauzAL5bgglNmZXwUEmbm3Q0ZNt2op8NmaHXnH/8V+pOlZDi3r2xud5jIGy+q7jbCkF1RoDxY
65BlwVUM5PmUMWcl9AInYIdK+QrlvTJu+Yb3vFskJiyn0sncqBTbWP7bSxUFsYf5ENeapFoQdPXB
4X/lxw1oPREOvNknGVczD+XzOlvX6/LNexzcs1ndJmCWOj908Dh5N25Cy0G6Edsk0mxxf3/zfrA7
OgKsnt2FePpAQ/QADSeqYYmnGZt8MGsqA0xyDYSYIXzXQvRjavXcjQLKpW+cI5uv0eljkYLC00Pi
Iz2g1+0R/mwuvpeRoDE+TuxoOT3Kyp+U1AY2oaxCN51TTKz5aKuygFud9nS1uE7T8JziNYOAHBPu
dYVVBIv5FxLTkJusJBcUzG7kEmptsQvdO1qEmpXisL0bhTiWWvgUGXSdc+sQeQrFRPxfpbjgO+s5
aQ+nWJ9dllaL63NCtRxPdkFJ40RP56X6b82E/KX9/UZS02X5ntr5fA+abxWMgqkEpc+gp1zPJt9A
6VC2aGMuxeXwwtyOsiwwi0mYcmwo5rVRlKrWCdc926J6qSbTiOHalNDeghf03/kBw20Vp5uFjkuc
JOPdDfZ651YlP/OZTAYKfSoD5vYUgUjjd5APOzJxgdNhH0V4rzbPEA3br5yDue/PimFaiRvhnz6a
fOagy1feC7SpugFrtk/EOcoLY2cQVwDIILw1qGJ2y3a4/iwroFXSuvEGY7VSnOk+VlCkHXO8fP+N
kMgFWWYh2n3NkvMwUTjj5VEOpd8xQj5G7MnHAhzLfK2fnITvvrvk9FGx1YxpLUgtJdiZClYyP4+g
uLmZLti/XDoZoi2sfFl9s7RQAXee4UXGJsOG87+h+ri4cEKh4fK8hku5wPy5jMWZRM0nKEbUjS5+
xIq2pyo8goBZFeCnpwK2NYvJmPdBDaBrXcKUePbe+xcE16G0GKeNyYhK1EMPHHQkJRNpJiQNBoHk
mpXUF5DICgOINWlJHn13tGJC0iUnvYrmaYf4lPQJ+vTTZ7kSmG2vDeu0yKWHMh2yBZ6bkheFhurX
KifWUEo1NEkksrTktYGytSaukCeoKJovx55deiyv0oLOznkibMrF6f+MR9CBaTB8JRg6jI3g/mvB
7OSHP3UP0JNafa/RMWADrb+1N8cRX1WNmv/naEk41Pil+Q0FyC8m1Hz3+fd7hhBCTIoiWM0YgOhs
nz6XF2qcQm4fvRMcLH+Oy05SxyTuYzsGbHG6Qyv2xTeqV6wjvEjCprTSNvltClZknIkv6DEVyjrG
07h2Mj/XAoSi0V6/B6dW2E2ay4OIn2AJi8hejDZNoyJFNi3yNOMw4M5Qzeq1SXJOvzD/f7m9eitg
cXL6kTH+iZ4VAE+CdaZYiMpJ2HcSaknu1sKEaQN6IadUQDxGbMaZX+IL0TpWB+hdB9HFTGCBCms7
jwev0610w5nis2b6sX4cpNAOAdznpY2h3jTAz4RKXjG+5SPy/57hSVR1IH9ZDnj1z0xAHLuciAPs
omIHSCbRvxNCVUgABRK3ibURWOa3QzMvCmbJkR3c6fGo+dg4tEkmA4FJTHF64YTPbqrlrb+dUbad
WJBrPLoMpc3eon0QAZ5GjOQfmUq37WpdzqrMB4El1e2EnoCh2NEUpt7LfIAFDdAqGjH1P7qBolsP
S/3EGyRsbdixDNypNw/0D8wR7suhWWd1WZpKs/tvFbcxy/R3qSAAJq3Ji7P3KnbVOYCYwExWVH+l
JBm71+USXI0/Dzl18YqZrSiJjFcYD/qRS/D3+fTeNdP/rUfII+rgvOGO6B6hJfm5fYhxBzD2v19x
bwpT2EeSNbTbCaNSALkzaq9bQXGGLb/b8h7nZp/v400NtwjNIr8GP07DMV0EA6Dg5RIdXi2UL5tj
HqCoxUZvzJ8A3kXTSSpJzMEWu5caDugnpFLa09DqGbamVfFmxGyHKCzR13O+jM279d1HxH0RXfGL
imPtKNoN7BmAkZq7bKtccwm3tF1WDmTqCn/ofNtHK1n7BlJ0cdgbxQzIhZK0/2/SmloJMZ1G7BMT
sjp4ILw+ZnlyqXqRuYlYg63UG1QpwInCrS61LsbSn2A/QPSFlB+UCovliY/s3cwpBiZdfIZumHNs
z+ndd/VFkxQU8N7I1MxdfEVWjMBiaTTIP+nTBgYj/cVvpgSb1UO+5TREIwcckrSaDbtEFv82n6Jo
IQenYWBs2Z26hvE+A2jzsdKGvEW/LlcZUtMHd5doH3NPbqRD0hfkI6ZiiZCA/7f+Uf0UcYYK9WKs
5aECkUOIovazIvPqlaR7RCMN7CgsfYcvldV4TYZ3YTrVs7a93qbwFEaiUedxCVI9xNSgY2uSCLsZ
baltkTaIZRJZPpXYdBjaUFb00tVc9Sdm033J4VqMGfGHlfutXjMAo7iGruzO7VbM9251WgJTIEM7
M7TviGekcwne0QO8J7TcJM8nh0IpH8PL1X77jTOwhPxaMdewAXREmC0hN77b7Hm3FmDgFhV73RGj
jZcREGGhEzfhWft9JKqphJQJsI2OYyrlZqAFOfIBMvFHdU8MgP/iwAX4u/JoaUERRHynrCjcJuNH
+s/2+nZSi5c6HnNW8Ynn55efRLKFNmJuy6E1fdswReSuXTgoHpjebcwrycSwYCFxywuZdgUmhMO2
5KkuRYF4uhAyAt/cxUgpztPChE/KTkhMQjwqu7W+dknnoaT/kxA5Zs+a+8jqIzh10na4yamFKCr8
IzKEEkzfELHA/+X+/qWCEdBkonqypCmqHLgqtz8fVC80f4lSEfGfzlXnBDfOYyBnJNQ5zpU8W0qh
Pnqo0aRqqFjAFfgCcjmWc21JpRL6UfwSdopB0Cxq2anEXjjeS7mO8Wuh43FR11Kq22VNPKl7O/yh
ujZSU8rujR18sFWP3Wgg8D0O7USrG110qXzKXRilDmLrPwjnLcDk4jsIm9LBVa3v+VlYBfs+BdAX
paRJJaLuM+UqZ7do3AVt20P8VMprvBa/ky5yyw5/SVjs9YskMwch009sw4oIzo3jsj9xIoG2Vqjr
/yL+4AlZzgA8/mSWzT5CFyje/HFje7KNOLcW6vnSr/15YVDTeNsW92KwBqC3P804gvu6jK+pQ2uN
eub0SJ8IPPpW4CZy92MPvnhfx1gDyL7FIjVnYqMhjsMp3ekkwigbYNdE4qWzWAdS7UyyVCv5fszw
yielc27ebbAzAAsOMJ0XJThsW62uZATjtGgWkNI92o/sl9sOnPc6AY2O1qMJuHIxkmq4Pf3RsJvy
JFSSAevhy6V93VN4azFilDrX/HknvbxJqVn5k0jcxkjNlRSb/vEjy7ULNNdARJGmXssKOvqr3zAV
vtC8wfv7EPnRd3Siu+8pfXdunII47DKOrIFpxJnHsrQwFByai6zGdd9idc72juklME3HJ5tiWgT5
xPuBU+Cg9xnWx7viqL/v6m5xqY8C4WrWsDDf7MpkEQrFIfxc7tRUTQ+GsGLoGka1uGkiWDT3I0+j
Ibidu0FbGsqR1zu7qJCg8+E6rGu2hhBt75xke04Q1HeA2QhDqlcxj4gCiK3CvHacfowaWDMuwCyM
L50aDoQ4ZYq81jPrV/HQpNh6oXkTZvwlzSvi7FGPkELDlOpCnyygAJOr6mS9EmvxBpQRiDFDD0QV
7Gafa8Zra9omexNfYbIM11GlF2qlU0LFCxoU3L2ZQHNkX3cYZIdzQpBX5TQ7nd+P2gVbtLOSQAFs
pDJZ30A6nAwPNAn/i2vfrzIZtM1OS5cgf66hk95by/mmUl2TQfzXjg8FiwueMUK1dohFBOt9qKN9
XOJBmVbEPh/e8cCJCN1wHZIntr23r2oI5O0P1XKoXyhLVsuQL6Oo1ne/DXi+D+kyTrkCudTTb91a
Ga4ouwHulkKaxp7xrHfchNLq6z3K2TrV3WGpptmpWZv5w/eT00kL+h3o6VfoT+H7WmCbZjh41iO2
DmORp0Iq5cAfcUh0Bg4vKAwoszXC+a2y6i+s+kSykGeg37DWGWZAQhEZdWwagSJ7ItyS1QZKquT7
pMkEstpUhgRJ7A3CTaiAumUwgRjN0ZO5jQDAboB+A+Q0Lzur5K1ua0Ejj+jPku8xABd43G08VF0+
vpVnYvbT1xwYUOwf0yIvFBaSUw/9i0v9JHwWImjBG3cMLm10MnGMdR8gx8TMnwMxojisPdp3QGYh
0SrML+R5TYlUc6poJCssHstDoIbC5OPpjpbUXhW1KBlaqRRGbM/E+Y46SMV3qZPvhDcFQNBq2fsi
lKZxl/xWy/1ftClSanfII+acjcpAGyTnb+se4cXzO7ks33SZ4RTaO1m8rjbcAXROoAF4m2cbCmjM
kxS7fzJEvFUi1EFnz6salYToQmzdNnot46dXDb9v9DToUGM4idOrpXl1Cgbq52ALxqzhdkrwBZeO
BVDWYn1kFt6oku4fOVAUqVahrHW0giAjBC+zlWVyHRD+NHxbPGNhQJ+D1kt3OOY4+xiDty8su8zD
3V6FX56VABaQj0GKE3bhvOa8AN4mClAD1iQxSWraUU0TO5Bfr1ejSQZKGMpBH6aHuUCPv5QnLY7k
3p9zxzqVcTTUJn6Ua/eX2ZNyG/x/nOwmMoQvdax40zHV8N6yQHndrQQ8wIjm/MkVG4Tch0xbGkG+
L7XKgW0Ks60pZVF3/ly3ibvcSil9SQSog8/jjjhfWvloXPpJSmrnY3BXBjhjl6ve3C6FvXuIFfOf
E3gFr//3InIEeHZ4eVb0AfD80to5a0hZDdwx2doI5WuitYGrFjqPE+xUmPog0ZG/syYrVaJ7sKf1
FNIgZO10ZbyjdemG3hkcyfly00KM7GS7SGmIm9KgKZtE47nHVneqJdb2WvTa4q8+JIDEElqMEqCX
KeL7Csur3JK1yq6v7CSBDCDsGsfvG8WRe8iHaF8DYEdQwlp+NQB1kHgbF19xUKvGJxKgTnbjxlRU
oN43UKjhqi3SE6jyHGIyo/Qpfy0xbyBv0eenAGC92KdKG1lP/skxeyAJ645diwrEVwRWff2dEj5+
TUfXCK+3uvjYf7lxK6TpfhIbU0ozh1CLqB8XAbwFjN5qoWmQ7T6qhJByvSoxkviSvhwSr1AY1ySS
a2sA7iEy7My0Kvlwl2IvhT0TAxVe7GUPuptN9rtkPuMEn/0IYm0U0LKs8Pnzg/SIvevZJaNSSPak
uKJROzLSmj30bAcmnKBU+92B0dFX1jNbOTpWHHG4HEFVBRxyKLgnx7gqkmrJAH67gs1qeMk1NFa4
k1FPhWlJHEfq2RGy/lTmk6Z2gYpkPjE09hchdf1DUVT1OvsjKnaJi44ntGlu1/NT89u8RUulNgHG
i0XHlous6cYpdEfiXiFBhb4qYtwguUiL2rtuqn/PZYGqZ56sp6oBWSDLYxNkdZpeHIFV22MP7oTs
qjQaEZ5EtdThCF4s5O/7MWA1WEkDcF1VG4PUIhB2zVXRMF41HKlKwyUuMVkpAfJhbLXMhzp4In+E
btpS0K6RoPFSFZlhJYpsJJvhZ5rCCSCmSq76+QA4DFAx5VRt1xWHII5A7G0pKTjM3FuC+/oc3SF3
X1L11zlXwbZSVQR4SworIbc3sMkzTtO/+qtErZbEUFtwjQHf/3DQEMyNwnLNkDaQiMTEcu9mDv3Q
qicU7rVqONH/UO4HuwNqrtQwktkI6tGbpB79VphN5AQ/rggDPEM6LSdNyowy0A1V6QjarjyLIXY1
VzaZ8GRZJ0i15vIKfpcR833nHDapTbHRFfcbibIaiNLBFrnZ98j1FWte9O6GBWDYaPf+GuQVHqbK
AvoSMcp+I6dMk6TXZAcf9z3TxNFW1/FGAOng7UotSAMTu4OhGIQaym7XT4eAvktF/7ubSlyEl6Dj
iEcT3DbTPPiiFsisvwTHR0dwX/nnr5mYF9wVDaAzrEKImLc/YTQyInQHitgr1mZERfyz12MGq3dP
bulgFRoCAPsmZbuDHytRb1Ol5qTIa0vC8Uibd/NqfP7nPH1Nn8Kr6NKdqcAHPrN7fn6nKsYFZb+S
7Xgj53mR5qhVXHtgNM8BtJWVdYfk+6F3z3HEqILblfMz+MqnTeCe2jdFCvhTI6odzd1K/GfPRSXP
uTKG8Jbsj+Wf8ycVI9DZyU3lDc6GOlAV+AUNhYa87xGdx6fhquMJNUSCDKKsF4eVsaZfiX+r/ztT
v6q/IuY8EPmThuMdNxgAnGuZpVnAjk3QUWODsfYhHBUK6PGD8r46OjvnfCMl8OjUjXfinKymn2S2
sHfGwnzQvarhI8PnxCQ3pRoxfGwZyP63nAyzxvAOSvsbWyr5gm40ijLDxvjwqUbjVL8pgdwvh3X+
TnyX8DggG+3GfzIpNECKg34gpHygetvLZyAnWpe4twSkppQFDm3S+3T+4OQkeAGnY0ED420FqE73
HlvZeGREUc4RtwZVzvxSGDC5GNn4s+sSNwmrMpKeFo2WayWalwomIJ75Yyg36YXEFg6hvT2la6Ul
+DdU4YUBxquMLwR2ftLu65obJa15vy2sEIJnVE3cRao2cr6IqTr9Z/Caa49vgZxHZRCdiRGm+6L/
d1jX3FS9iI/ELTJxJgZMK/ioQOGVAZj7PjWxYgs/+GYmHc3+E5sFMi3XCZ8bn5q5qtiBpfQX/jz0
njws0aDHo0qDrmVATuXikKsXPesvFuhpFEguijnGMnM8CaRRn7yBywOZjP+kC6sEU6GWRKLfbRtr
Q8NRMmh3PrTveSDk+2oecSR2wwj7elp6aSXsV66jBduS1n9PO9xiv8SAQrCOkYXPqaXzxkvJn1xg
ACD4k4mfbHyQPA0YBsFw7tGS60fGNHP6qwQhrut+NQuzQ2xdOLVeDfstaqqb57HFV0VgBWYS8cMf
YYRDHzTrUlMUDv+OCS/HGQQrBb0W2BnEZ7/p1k3VcHWe+mD68KYimmTLf+t5T5rJNm/K5ufquXbg
BNc78XinZGK2l+aWH6eMLQHsnbXjXl5Jx1F1JoXVzWUrqHayFttlcS5KdcdoaxepFfm5G/LV1s5u
e1tOkvacq/8AehUi6OpKDV3vQ52cJQtSFwEORsJRV2vLi7Q7XEdmmN7WBPot9ZyiZwr4LXVSQ0Xe
EUg8cEGa1VSgc+/G5pc5mqYzTU+7OwNv0a/jvtHBWBuv4gdYuUVTXlsJ2/t0toCvGzn7u3MgqACb
4II47x0NVRoi3MiYVISKBialzLnThFo2EcYXAbELOOlJRTQIynLon7UYsaq4m0x5ViM8C9EoRNtQ
rjqlp66vi8m7amuDSDabXpChgB+lFIi3/TLapTZFi5/W+SQntqMziFntVlF2MPhfaPX+cGICnQfe
1GLFine+2Z9VM3093h/cMKjb4EPSu2MymxfQ3xt9gN4cs+uPy75tq+ry6ref+vV6d5PP8wtgpsRQ
EyrxtKcDoUdhVxG6XB3QG/uObg2uhAFwTBuuQwQIo78JwHlJW2MtqicQ5Zfs0CtGC6GmnAUEGrm9
YP9HswDhpQOqUY/Y9+ZPA65k1kcbJN++z8X2sC1xaAGKAzoMgmZr1PDI1iLhb4ZwBXnme58DmtZO
I4QAtr/zhxPl3WXjzZyvp0hYg9wMIB+D7KZuJxJ446iSB+a3YwaU6uKbJuV7RJlv0CG6zWnNrGlk
igw+gUV4qwoMqeUJruMQowSOSFuYfm5Ef/+nPDS8dQ3440SeiASi4RSBkD5HwA75/m5MQkBoN17r
WF/Rlp8l/Xykpgh+oKKMgV9V2xD9aHmyeB77Ii5NvZLUz+2M3+c3VbdBlmH6LtzPuwQ6xr8dmROy
r87yX6rMQdNyxGL0G+zFAu1szq2iVV+XVO6UZ7qI25bTiC4oAJJ3AbrlOoL3yKcsGVWKjG8DtNS+
qN+ma5xxW09vKZst6N6994fwFEhZg4iT69hXwGTO7vZe5FK43CK7ewFgFtLt+adm6MxcCZj26UCC
aeUSQ6V9dq9L1tB6lbOpcY+Rg+vLttRZdBe/8Dtw3KXUKCsjN6fK30f2DJmkhEavTSrg/EmGQ2oc
B0mKdEKwB4+XMUrpMKbegcxM3PhSLpP+gVLXsIEtQQ40s5FPMuONRC6YYgZlFAlGDlzXWPYHkpvu
mwW6B7zGOoo4Ye01lEn8vL8WjJU+12b7shE70gB5fmNQaZm0X+rWBro4e1YOpgcwf4fcfM4KOzon
wTqvo1RxSBcBOwMxH85T8osE4nmpLLNodDMRP+MVAFWUmFEViiPi35oJR0E8FU7BVioN9so24uQm
JiisY39LcR7KSnPcUDlAjp6BOTsPsqxE67vVyqL13X2IVVHDqkIRgC50YuhbZ5WvQznlPwuDnjEb
VIfN9STK9EcjeciIyYeMoWWfwSajb9uXH8z8EOpVZmMSO2NCyxx/WINP7/EViW7aHszftEkqQQlf
pCIzXr0jbVBTerjn0hIJ5N1/RO0ee0npE/tqSlepnVclDQtpyGUVfBQvhd1BA+9na/TmNqnP3po3
B0k8FrrNSIDOtT9hHEFOlrhTz/PxGCvPg5tjMbZduUoMACWQNdgJL2RPKh5ue5vCeYnIgbMPZVZR
Ulzvr3goa8T1jY7wyyU/15+b9emvC9Mv0/wh446eLjXuApACVU5uM9sB0ZvYA1M4jUj1+TYUwmiE
8PMRmNxp4vlX24bemB52p63Llzls+8hj1zHY8l/7KoLufNz3EFVsjLckBFtScgemK+cCdB2m/KpM
sdwu7B+SWoLAejni2gyy7MEOs5bf4RwB3eFFuuRFYlct9SBMtgq+CJ6z6G1Wxwn3wjbkn9sNLs2j
7aczk3MwtcPXDb+a/IKOv7DpILAZwkwuor+tZeCUMJYehicot+Fz6R/FrAjq05bnZ+FW9iwf/wHD
obdszrTwbK3yLuHqWHx/rDZLRNCeYW5h/zlejaJwHAXHfH53/q4CCy4zQXTl+1daKnasoQZe/ZdT
3YdJ6iBEONdiVwOmXmGwBgl4uXYnWkjn2zXbgAMp3PXjEoRQ+ngFuqgO6wjHsqvi1YViinHYTgs8
uk05f5TThBe8JNjQSSSshb7GzD8/9Q+uMoNjPxb/UeDCRI7YIWsSWSwuV3I/d4DfEUPLGfpYmwti
L5JeD718eDYhgjYZPQFRXZLpeboXEPqzXOm59rDPT/sBHqNq9QxnH5TDgkjqqg86Za72pCy8D85K
hr0YsljDUiQkxfVoS2Qc0E66dCB28WZ92Jh4/ei45vviv/b1ckj/nm1zDDisYF16iDSBadbHzH2Z
vgrzjxbht3uJKjQl5AC9FyXFJMJ1ubC3b6iaudeTll4UzBYvbxwiCy8zCEgXq5d2dSqtfr1D5z2v
9EN8+3itBCROBp0KnSYf01i0v9TSxqnZP0WrXdY0jYA5pWVcOc6JYnRfU2badC8Gp61SzZUJsySl
eEKlELp4Kc1DREHEkzjcGKIvMcDZQzRgQaPf2uZm+XdLyraPadPa9ujC0zp+iaU+apRBd6vncY+R
zmuFU6Q0IgYGPARBZis0HrrgPJVPsj7hgU29CCCgKYuhZ0SUDX21rFkwPl/OWeYeKGTne0kHe3ye
0X4hpAsnK/9JYF1LHM3tr0Wd77TzKkltzHMyTQojn7eTQeqkVXJCrhaui0iHvk2u4TmTRCufsgQ5
ukfVGLueav/SolbE7SYSsRf6nm0t2PgzHF9BFVyDAZ+FaGClWZxQoJowoWPonv4ZX7sNGL1g5IFr
Ny/ij+I8iCzRzchEnKJ2L9hxXWONnnLsu4bo7ir6gclcbcLKDW418gBGQQnCGRJr7LNZJXq92uU7
27UEueXOhjUtruIEtsqvE1XozVfHolrCYx2MaF3cCvIX8NQ07WMEnUIEjPMO00CVIfx+FwLYWasv
YAVbgjgEEDq4OW6SZannPs2oBTm7US7oV2nanfjXv4PEy6Eo1pzDIhC1dcEhaO1DkLXt9F7Fzk5w
PxY5ueCMjSmFNrNw3gyyVg7L8XjtXpkTEkAVjpp2NK4R0v8SMuyxdxyohA4NEy4rXwRzwKgBZ2IN
ALJ8YrfqB8TrsJczodCmyG00/a77Q4Mxqo66Wr5lAnukJM+qwB2LXoHXZsvQ3qtSUvoEvFE9m5/l
MuUFE1yJcUx7eV2acUg2Ybg87vN+dkuXQ4sODti2isDIE9JxfVnebb7RJzRn/qLe/Xur1/8nfpAD
D4XKPlAZ/0nKzKYR3Ls7nVFbsGa04bp2D2P2ZIFsevkhMy+4/W1KLi57xG+PoCzjQYHagVxklP1s
V2YHF4ykQifgwQYYt+XGkaADH3bPQ6gvHgPGqrdVieeNkQMDzMBGeEFmdTi1niW1Vnb6YI1LORpS
gxdF2fUBavR3ptehXVIfsrPJ0Y8rGR1rKxmdNnf7g5F9PzdVhpb4PiMfzd/sWxbdTVPuKLLkChvz
xjbAVbJaQ09fY0dFjAnkDzdebT+bVu0MrSaLSIh64DqKCfH/D3Zi7exFjP2b/x75pws1a6zYwYoN
FCzzIcLZ7+Oic+hg8BdHFVo1IaME8TghXpdqkqgccz7IMa8chNEKMKe+8it0zd511iCLKYTsPxa8
T2Vp1q74ccmTNeXSmpzZINBrBH2DjjniHbfUeXhIsbY9HVuZVFVvNC6XmhPT9g8v/aFUjINInJrr
Hyj4y+Y6g0kvnRrojFIjJuZC9yskaKHd1UCuIT0FUFfDh6/GeF9WdkzcbVl2P9xHjPDPG9uYS957
tcTP10qeFpqt0zLj9W1cVkXcf/89W6U7ZT0kccS3ccNnzf0bmp3oy/PQ52IdwCa7X9FtvP1KhOgn
PoNX9pC30XcsFZtw/gXcCTCntGRJT+oLT30NgxJAfp0ImS//bpSqXb5w8D0tHeD7SmxbZr/tp3Oi
j5gqYL/xIIjLHn0G4BOZPtrWxB+t4C0QPd9FBBBVrE/t+me0/UfKXxQ74ogun/9TUJk+lTZgWnie
asRlWgRkRs6/yq6lUL3FK41E09//6o9637Wo2HDAONAVX4AIW3A0SS7J/lidABmFcCLrV+ioLqK5
rMI9eaLBx0VYa1oKnK7R+CUQI7/aYjxnE1TlpAhUtihe0Vo1kM1gakbocZKAKF0mNgrIrSRsL9p4
p01AG8N8gBVzHhgdrQyIDdMCam5ZQuaDvlUKMjX0VArEGCzzQ7u2tgeyq2tkZlJKYntXLpQfh3pX
wIfslMuaJCG+AUfWuHTYBbwPdPbPxG1RFI6BmpXNOlsXR/VGiUw9bXKHXyfmUdw2ihD1H0bMGyqs
ihfY3/sxr0MMcf3dtgZM36Orc8DWQkKXe8U84oYNAdLlbhoDO/xQgx3eVtsRJn5XbFtTb1Ig+fxf
5ghnvonpAdTGzt3LYsHMUU1KAYonW7Lg93NES9X6BxtxU39vR9PS6wdsqQqSOYsgLy5ZMQEio1NF
0rHtP6s3dbrqJuLRLJgK5gUJF31ZAz7Bt8uRA3x6+Q0ISjER0Z6YA3hR147ZZ5px3pLCquAPRJHv
F3yOJhZCRwCY0uDDEUrhtKbRA1ClCBUS0fJ+X1EQFFTXbj/4l2Nwirq+Cpq6G3loWZtfW9q18yod
W6yRQPmpOSr+7/BpVcMjRRwo8Wf29Cxx4769XmG/b5VfLd6Wl5oXyYKxMVdBLTLn+L2/tVekLKPW
YlwLibqHfpU7QGc3LI3y8WNq6ZTdavkC4rjCO0YB6ArZ29hgraDymJ8Zszpbwbm3rp9GuY+HO9Vk
USFQqVwU1PtPtuvu6x3+OzLBQC45uD8mQ+lnlrHV8SRqnqjBthDVPZNxQ1hcDWBXQPV+9MlxvV8i
s576mKbLte4UQ09onYuDXeLyTXy4shLy4awpXzzxN5sWDutoK/Uw6Z2w7Xabo9SRqwoayTSGvzWt
foftK96DqMVFZQ//2LJTo3A1vOvBTUCfazP1IpEU3dng9DaUAoUOMYZlamJkxptywjmRK9cRgyOb
nmfoUygIGr3cio42nNUCo7nNlANJBpwRbTMlfbzxJCdDzzvEg/OcpXz+RE/1MiU2Y/JtcftWNEIW
8ctY+GRXIwVte/K/oqZ3SmzOM64DSD1OcL1WGO4h73rHhQ4xU5WprF6TCBOVnv0vPCJOYfgskX9a
nqwh8xXfMR59GeAtCWgYcYvXEirWI28nb++WRAkXlOBrVr082oTrBAfn6XJnFydgcY7BbD5+iSx5
MM21pQ4G/xgSshkNGQuSgsCtuEiV5rz6tyDHKv64RiQGu6YNmjCV9KhbSSyiH6w08RTOCAzOmGpT
nVMaoq2C0xKw+K17Ppx2wYWigh8c1IvvtUNrJi8gaOF5tqSr8neNfoOeQ2RAR5njsZ7LsohyqZuq
hkRMLL1hOqGuxbq4R4JX9PU5QV9Vl8s2vvwCMgQmmdUdylPhORm7gkzRI5CWS2X9YWHbX4GsQJ7j
yCx6dEpKuuHWjueAHFHpWDHvxlsnu9m9tfAtg/AOsFjaSg+tPraC7yx0rznM1GXZko+YdA5kEHFs
GKSaWwsdt6gf//ndZItMBC2xULtQwESJfJc8+QlQ+oAlk8QneQ/9gpd7pKvhBepRhHlzFPgYHH9G
rUVTX/946zNZiUA278GTCKul3dEZQDMXEFWMi1OCQwN7tJK+H1au0UUm41W0Dbvnhd5wpGuYRplf
GyFqhaf856LYhKik3Dfsx6eyukawnXbdYzy1vtrDrfjJZEzjrnyg5lnQBjJG0ZKSwpjmN1IAtxhN
9+jMcVmlsiCiN94XreSQ6YbmIEAmAjqhOVT2ogFA0Rm1XP6y74gBhEpRwL2eLlUiVK11QnteJo/k
ixa69wkjBN2LkNVZvT6gR53jkMi878KKrR2ZJp1RIw3+tTFp127+LiWpBKtZWuFQ6h8jXm49fVrp
jKlPFjBqbIVz3qd0Sxp3aW1FSKNxbfbbeE4sF0N2Ea4vvmvBWnbkbIY9Per4HCAGqJgH2EsvSf+D
tTOB1MLfUamlkoZVYOJGs7TdTRWwVZlP4SSLq1ZoeT3aELLW8+y1g6ta5mM0n8Ko/vtOnUgF+AKS
v9S/nu72MDg3gIcznW/VE3dePdbbsOFk/bFRXawJoqRpqQnZV+xfTmcNAhYAp5uDsCtt1pf1i7nh
RssIQU1t3AtGGF0lr13Fl8McGv3/GLFSioeLf8JEgvkKa4uJ8XKYpI7yGkJYA4Y9rSId9eS02JZ+
I2jHvXtf0MA7KcPYnaEWBdPh/sp2C1/rS8CgdiFqM3fWBKFYBqq1g4/V45B2x3w9i2E2ujTLdQ2S
pbUCfm0lSefoYNoMnG0HozExOh0ZmgxedtVO3iaz/ULqd/m7dHGwiGZUUs+Qk4f6+xWiZOnyk645
lvI27H3SdZPQ5DXTk0AA0S93R0GJLEQXkuCGZ59RAmsgIT84+zGRm0SFHt/6Ny7x55N4Wefr0Xkb
Tgao+YyZHEyD4ZhaZywFd48KCUYit5BZFfZKgTFdHuUS/lbxxQjADd5oOn5XU4dWe8QjpNJ08RuF
9YGKiZ1qGaZUcX+h+GUtqdU2pwP6qnVtmmNqhO+IU28NymEFDr++bp6MKNBXW++Pdh9bqg+cESQy
9LesnQqlojSBXkYD7gQyfJE1I2QUIcHPVK9GpEQMW8eRqnJif4hi0th1vkLyU6+eL+E8yuX61y89
UYyivjMHv7jr4Cca+cB9w/BNJ2YLuFk4q6DREzS2s5fFZGNoYDIbUeHC9KM+LEn2NRXQ2z3KlqIK
PzGJpdDfxOcVJ0+exI6M7l8kWHeSFRiDSko2uFy3chprm1WWvymmSnzs/rmfBHPtiwb8ZDnuLy7N
5oMYsNs5ld7p4qxSvZ5E3FjTyEvWSQ8uqjwldybW7WbJ65yjyXf8dUm7JdpV/l5QRpst+Ui8/q6J
6OgRkZsWLEktkTgKropx/7pyB2k+OYZ78X4EMVwbhNg0ojyt2hB6kb6zteTBJbZECKu3HRUdqynY
mUJ7H4t5qWYYYMDnxfR1X19T4KDkzCD11J6zS27MnxfI2v5aI3gxnpc/6AnAevBTFKnOdtwsxp+d
K+d/AVFgoCzpO3Y9ebO2FSdGb0Y2HGU5UJT3uiDFPoEw9v1PQQeEGp4+w7I2gcgcP6ZRpIL0poIE
gHGO72A8AWhE+c1OE8PR9KPRmeeqw25yPIUSyw/j7NuK9Yz0JykPQfeVhLcwR7LbVItpFykxt+9t
8iLPt7/wir4/bm2NGZoOq2jvs9p7NveizpBAARCwoe9VUW9SPz5LSxcj4+gyGc+CuO0297VfV0Hk
/Qz5BOV65cZCP1WvrgX0toROiTcCnDZNNKznWwfsaKSaKhC4Sy7aHpwfpG21gkAxOUcSG5LcxUou
vDuncLLIg0onTc7WK3/4BkvtU2oFuwawI2FYGXNcEjbdMyYIEnzrqE8D37FB7+kQQfDoVR86biLn
YQij99Y0ZOI/N33X+Es7N9aGvLSlZdlyWwvt8IvGPdahs57wM3MDL7zk2Sbdky0vmAUpyQ3mjDdT
+CQ/3cBjg3FBvvwyq2QsW977EBL4tqefjXIG6XhjS0P/JDqaDgslbznFxyg3f8MBrqjhOYOYkObM
tl6XP8kzy3TWchqCYs+Gbv9ES/sld03NzFPiuIScPS+BwXqP4qcCS2Dqer1kHzm+tf9gcXHHZoyO
RdMtL50FrKuDx7ZAhsjqX1c5Rodz00iF2WeA4B0MeB7btPzdzRizKD971SogO3xBlbu863wFb4cn
GLkilk604Z7YOMMHwLnO0wCmgXn3a1NebgfxgGNP4t33n414cnRpmt7pfMkgzNpSDQcQURm6Xde4
H8SjMw2sypMLcyitl2fOT88MIvMYY+oEHVANsd5YqiBV1+f32B9NhicSyHv0u0k8t/SBLu4m+Qro
IxbjBkE1GMdRHnTkO6DWINqeYTNL6s0hrN0Xo7uuJ+cjnFaTWpx2qeqgU7KIHXHEu3uX1lJ1mL8Z
zeYhgnsgfmHG7pXW4wnk1sGWv2aRpamWyLyVGYbpQMwcCAEXkxVL0k80e9ylbl0FrKo5AWFcLFdD
g/KZlA2/NMX93+joK2AorN6HL4LK2UlDUlh+wlnN/M8aX9G4E37NzJ+qUXupZNn4OW0W6NeHnYWC
1HBqVJot79DAIgEKveawKYmp72Sgw3VWThMHgy/4ZrMN2OxtRMtLu9/LVkvEEDeyBd5Vxdv1bO93
Df4ltpw/GgZqfQM8SD6Tbj+zB0zjsBuIGTh3bDVXWFnfmfLiIa4aArmJrKGuzct9pNISLDuwd6nj
JLK0rpzBB2yCMuivr1EJ2c8uKOxl0kMaUQCgFjsOxhF+hIO5OjrIBgq8n5ohgCpUdYiLFXJJX53n
wlk6JCvizzCqZQ6zqjPAIzM3B1CLfGPE6JSFJ9R7Z9ETay6lg9eYkVPaxi2N8vbnTJDJTVnf+k4t
3+OoLOEj91mVLMd+sBbMrMPecNSjA3OW3bba7pNZgZxfibTmLh5UbFy5QGZcQOg4Vg5PsWtm6aK9
ncuSis+32bvn7VWrDIJvX+EI3iXbbqqFg8L9ar+jNmG5E9M4PlAHEChaQV5GLHP/sm1q8Gyvw5nC
ohh9kW9TjV8ypKVYSMe10fFgw8TPpRv3EZGeW99gmVm1AuRUpQYjLMFadgptMIjp1X31LNJKb40l
WQT3UNHdmcAia9gMfgas9x1XYBsvCIIATvsrhJZJswnY2hSCEENKyawfzWMI6X8MAc16quwcuy0Y
T9zzg8KrSrAiLRmNhKSwYD756auonmVZvZWAmOx9WbMKEOcjHW/P3fY+AsbZ9oXDJOHN88dqRSs/
kbk8CsazA002WE6HuAuTsZUXMMVV0DFnnh3uNE/3EUjHnv3b3Lsld7PHCqwXBKEhj8ge7UZJ5LY+
j8z3LJIUo4KJdgjfGTXqCIaMUh8QLLnDPckE9rQTlvWe94326SOPnLaomekflI8A5jszvDy8/H6O
OHZeH9UXCe+r+z4rOIYL9LM+dKj6/ZRFX9hQRGFRqIMqtcoF5/TdNATJGmLNEZtsLqESfw+WlCjR
XIA8FFt0NvAZXBnPupla6YUBVn8+Gky1AAh/rGwAWDT9onTyhLjScxmUE/npzHntT1a5KDt16Mv4
U6CWpoaF6rTjlzZkLm4uFhwZD0DidZURnogkgG1qTw4sRpGJfZ4i+S9ETBd5UPqaSp3fYFXL8BTk
mPCKgpx7Ek+MdvW5WgA8DueadYbsrdGwNcCLEoszvZ1Wg3nyiPMKeCdWSJmJKBDsE6NAgq/JYnuj
wNmRhZbTKhRicNC16KuECVK3kYY5jfNv15uuDVmnQYrCHGM1FEqSC3F1IPDCfjW/cnCj/O5Vy5v7
GTMunUw2395XJ0XNYjKcwScbd3XJ96+8j/Lb+ADg2zVt0iAWgYsPUMKhMXT9E82t//cXXbK7jPV2
VYCOSn1R3scn9XHn3c+w/nrgy4kBhYn3pu9tDcGmHTanrOCy9lg1A+dY0g6ZTrPncXyjZe/nfdi2
jvANT0KbhvfR4Zrnf3vLJId+J8GpPL0qyKh2h7Hxccqvj9mTun29MRO7auArrhxG6/GlzGo8hNAj
iakD1a5DHYUuymyWnva2TeSqNr89s/wUMVZhSqho66d/bQaQgOEO3e2U+wSzB+WfaM/HbPxI9Ngg
HND5oHlLkqNbh+orGfQ57BK5qTlRzjV62urr4j0swMVXTdpn4o4u//khp8iC4Kn+71YyzaS26Sr9
AT4M5gNqaaQOHG14YLFaN1yMM1eLNfltuZz8We+5e/WaShNyAlfkZF2rApqbt2ikde4EZlKBOp5E
4om+PB81PfKzVFn2JHWKPmgQU0D0pc6DSNNbdkEy2GU2BAx5vq5OUcG4nn4jY9xbPkkmAKVC9RKD
BmuBVQz+TbKq8jzZz1Yln7Bii75ApG2zRBDh6L4d8Geau2Gf/bV1/NtMIzfzaJ1EoxtdmDZNDhA6
vYqvKeJEEgqs48LKRiuXk7ptxkopezAIft/oX2ws1xa/wwrI1SnXSExaZfoL+rlIIP0W6/Z8ztH3
tE1afbkmjEjk66Xtl/rHLOf0bp+ehfktCNgmQZqgv82yMG+BmglNC/FLb/umQacHIJ+SV0PuNvcb
e0ezvAiHN9NxjmHq28hJ+EtfTusdCoFMcVAqYrl74/mCcyTVHFmXF+QTt4FZzSNlonsxd08+MA1d
dzpQpsN+GsjrncNuREGBf0PbxN22mPucLlf2VgLdL5DW62TOuGUcNC3OjT8dsgnkBT0zjhcqJ3bR
atVNycjT/wJSpaphzNTpX5Iain3k5YPluP8j0cZdCaw4/zO4uoypVOQkhDLG35FsWhHITfaW37gt
0BNpeApstKmeJ13Br2dErbIdfPw8gO5YdiSh//2xxPWyKzZkJksTvjyb7z+NrtoqnaCy9hU3/HGw
SMAVTLeewr4wScq20qq/uTlUM4+tHoltp+0spQ/9ZkNdo6i0pEK0PoqSityGcn432gzyV3IsRhui
C4UMR69QBgxAI6jfqQuyT7x+E9rlcwurxbf7JpbIPRu2FgCOfaMp2Hol6YaScqemHk+tFJ4C/vZT
YFoZ7HIbSq7bFkJXOvu6roSOkUCyvkGenF0Ru1kTxQiYZT/tFWTr8YKquXNfXFNfmCWwnPx5FXyW
8apS8JdFJmMOQCJAgueT8gGEBJZWRQtONnG5sRVroFd5/HU95Vhl0cmugqiJkgsHE2qJz7R6xqKV
myEN2CqIlSwhbGZqd6YrW8GnMBIA18xjXcjtnTV3dZzxmN7nF9MRWbEpcPX9KJ/BUuSYUx3xm3a7
OOGFsSrMaQ9sWSCNUkHN2UH2hzgmTMaqORpCyrL8tZ1QgHUa9GVcOV+r/6Y6omJ9y4r2h/5YkpwT
l40MO3vERw3WUBydvYjkmIWSDExs9LrlgFYmU8t4E36N60q0jyyUiIo1SU66nEJYZaxD+OKRYBEn
SuzpvTjMQv+FmQJhgaEPa9nLJ7HX9jFngKb+14C4PvhqSAZmR+MXq336l/aEkkLd+BJNRdXeOHSi
AhK1D6uWbwrWjmkLNGjt45rXxpR0LcBrA7SPlXGImpR0u9FaZa2PRQMOOnuLmYaqnZjsmR6j+jhd
gnTA8+p96jmbBJiH6Va39BoXYKGXNVmPLrSlDUIqZiQC/aG8ZFXl5199DVRg3gDF2J32e1lcjixK
z7gOK6yyyqSCRGVmGpBkDLHIqDdz1m9c4iOpoP7JVB/iz79PqgUm4HianUCyYPgQWQLKUqyneTRP
/As1TZzIWQBItVgAmCnyIuGfpIhNiR684mzkHNwA9GnyPlUrB9r11hfjwOKQzgesvrnBgO3fijji
0IzB4x5cp6xZRY6Ewarcela+IPZZvdOgVFJ58EK3XHz+BWVCw0Cxg84xJ8UJtMcwz83b5VrC7iOx
HSfoxqEJ1LxaMBvnWsmwLxy4qIjVyEiKugnLGb2HLoHk7ojD0E6ApE59CU9tPBvqtAFusMGvsYSH
4+oWE7amEEDxZbjxFN+cTuHsWD6VdioOrlFcTGIIuIojxp94TZUjpkYGJ5+FlXb+Ekk58njjkCUt
eVg9JipnOc9K6bKzL11dpwGHb0t1GHbzFNugy0P3gKIsd0Giy3ecvnHp1zwCO/rlvVAriIdYezvg
hBPdInrozeboZoHZ2vET4J78Chfabi1MOX1FRNSirQLyeLqjfIfGKpz6fxjSsPScn3ZBiTbD38Ar
ghart7X/zR6CPTTHxXD811qeDCcdh6hictS9JuOetPfTy3ARH8fXcRI4BHo4T8YfvlOxOfzCn1ap
pGlpXY2QfXboe3nMy5o5418Ub5RMfBd6w10G5cW2vQ/LrNVQIke0JQvbcCeJxxjcfGrQCUvr6BQB
6YFPRHm0L8sTkmmtx8AHhc6ukHKUPF/P1AeE7HR1uJqNfLKImUuaUgcxSZIdk6GHG6IpF/faEaS8
vjdH+X1zrhM0L7hYZJ4GEw/O0Mk9oYGNpF081Mufy0Vehzyj4rSpeYzY6gHCv75C57ToI/QSb1Il
u5IwXjq9guMjGHUgjIIX+gXq/IkB3MjPnqBCi92nEPcrjG70OkdAOQ98u0nJnZllaPI362zhf6e4
4YLOPTX2feJN0um8J91yhKUstPi/zALaQL83tmsEmZaS9ZoyfKQyg6IEN+PKNNG3o6qymrr7KU6q
9B7Qad8dqfJam6CIXnHBYJlkCWE7FaOPRXk00n4JtutkcoQql3xWLAhhzPoaywVHhMFN1vrXOjFF
jGr9d6U4dLpGVKkN3vglkewvBke61nrMjNBZfYPJ3Np8D3j9sFwuDDmBQV1zFiOdVNbBSoCEQwqd
5z9ozT9Z3jxS3pNGa75xVo9cQhrcwe4rIWKTXzlifcPo+NoBQelbJu8Rkt4re/5dUzYkEphMWNvo
ye08Rh7qJsX2hANm8c4ruyQvh+jDMCCweCLAquls/s/OV62PaazgQXymxZ39D/ZETq4cFF29CDTk
XiG+7N09gC0D/lQnsko5Zw4I5L5UuKP5gCh9WD0bDeSLnn/LOtiQdK0LIq60i6pnX+G70BiGRD2t
BQCPjNWIaXyaOcFRyXwFffbCf8rjWKot6o8+h6e+pOjofB1MZDJyjciwmQFoy59J+alCS58U7L/t
tX+Hx1tSN68TrgMt4ufJQyFp6nA6TPOyzCiJlNInBzd5Uttn/S0pCqknM65jOo+Q7Dj9/aWcu/a1
5f9pTd4mO4w9J2qNLq8QXlpaTfMGFKDodPzsFw+q3B4jrQ7+zOx2RQP2+9/hpK/WMu1QjCfedhX2
cjYv9Gmsm+ZLonb/D4T+xmgffeLLrpQrPd5rHMc99839YmOLtq1TdSRyHIpGQh5zLEo5pbbAWSIY
rjy14qNPWK1wf28jD460nR6lfcLtmzubSMmTyWQeiUEAblLujXAzEzCwKgPW3MwL4Iwvv/om9BPz
f2gL8RLgV2b84OLTlx/hxBHtWtH8RjqEyCpqIrCrWPQDyA2+BJqHpXCsXaeK1SVpio4S8cgWY9JA
zzzFhPhyWJ9XoHmGCD+Wg23EzPN4oukQcCbIt9ZJY/mb2m258+i6L4wxFvHPKQf9cVi7pFPkHDy6
W9dO7AdZsk5RgytDPnkJnuCQXn41VDIxdr90rzrjKZE5m9VTHpP6Kc+XW3PQ4NHdDyy7sKCFNiHR
QnxdaC9nf9+9psZU0qSmDIceKH/8Mg0AWpY/7pCQs43z8OlSeAKLamAb0e5SKNNyhmwXBU8jjFyb
6S351nKTokVLVqOcG1n2ftaYKyq1pQE29/tzgJxsOb2YK6GjeQKxzPOC3valpLEhVrEflmseyYj3
v1WRF84RDyLHu8lrwGUhiLgvmfdG3nez2l9r9gqiuH4FQen/n2pcQCymWB/639xa/P97ARwzx9rt
Fl9teRygcJPegcamypxXBbapS0yRHCNobw9k4DW42y0hTqME3JE/7NXinb9XaBLFJI0NgWfcyEOa
+EveSQn4buWmf1Tw8f4RqJFEUk6GisNed/ZOPVV655r89Y9LjlkLU9Lu8A45cMsHWAqDxn/rB0Co
jp+5Pm6qRo2Htc53Gbtj/wNLXgJm/myguBWKKIv79+TikuYob69r5XcY3i7+rTweRKhIXZyI1Kvl
EkHt6iwvHpWARWhYeTvudRB+A2F1DMn8vkZ/IJt2ZbXeI06+vNZWKA59bhH49Td3k7Kr03ch+L/R
WnaOnbe295OgLlJsnJmL3mrBFTL3M3qu0Ac3bz9oQ6QFp3YGbTjYEXTPhbbjGprvurnbZ8nAd3wF
+OIS0r6ZEfQBO/GFxBHvwkLTEmcfItdxfb5dhtCMsH4XVhVFQicGT4GRHMLOMXOddJiHCquF9L/P
exylzemmQdy9nqkxQRFlo7aqM9d1DBnFGDYjqKpHA+iAgi7QEwENqJ4mzd18QM+wVVEbgzrE1Ng6
IVl9GxriMPgzU1keKD2idof325H5UyjjUduAFzDNbJMwqMzJ+dqoHLTGrmvvO87r0PgdLeo1VwAZ
3Uoq+MixUZAt8k0LVYEADhbl2AbdEQSknjmB8jM9VxJSfJlcst+n23evuPhw+GcV4dG2omoMhHMJ
LRteES3uyhXnmKF+TChMlisKHmYWHLccFiT+dQJ8LBQ2h18nCQChuFAo9mzibCK1TSXXajVqhWRg
+CaPesElkIQwgVRGWqPtPUGEo1/fxqc8btt6YMteMtfgK6NC6qBRJ8VA47dlsHDf0/c0t1rpFEX9
AE74tXkITdRAaqB1TmkkGF1NJ20B0Vxve6s6jjWVRjD1TukCgLfp5gTLDAnEq9oKu0Ri1sg5DwQG
gyb7c6BgORtTUIFPnjbRGNSngNtQqKwZgUykycEmb1IZCBw86cF70OZ1Qw7C6rG9+SnL8tYl0q19
PSuAzFG0Kpl+e4X/akHdWuvtZtneN4MuSKqHafwUMX5ONBTnjC6EnlLF1Z/zNgKhvs4/pqyQ1Fb0
DKam3FXs0PHaUy/3b5IpNTQ8hpEkZdL+XqXvgzwa2AlXlCtpS+HIME9zxC11Q1R7MYAyh3PTNXrb
Gb2ulmLHHthcgsurEx6ShazXDk+E7CdsfNuaoYebtmMXh/K3I96LkKS9oLQXwKkWMjBe7/snWZ3T
JxZ6UUWZKwg2+KjDwji7REaLsrTZwiIEpunN/rnrF/zriXHpNkrC2ZVqWETaqpji01bD90jWKiIS
B4epwjGbNaxyWy+auHV59SL6kpCvOsB39DAl9UB5AM2i5Gi5YfN86Yre2XO2SqxX2z5V+s7byB0H
xAkNGA3mJz6R8+jyEE9eepAJ55suWyVVxNLqriOl0hGKNw8BIJiNC8o0HQ51Z2tX+wK4OapDGN/R
Ss4GKtJY2ykd5fiDm7Q/mJm16+6kXr+HDYn1X2YkiYqzgtUMVca3y3BH5/c864d0VU2vG6NJfKXt
tXxtgzIcwevaVnDvLvDgXnNMissiP/llkd4QVW9kscSHbBPafyHfqWa65vxFRBvYk+N79iLx175T
o68j5BTCfsnDV1IkCG01NYJ8SnmMPx2q3p/YdqTxootdHlWG2qU3vpp39StI5CjcS6oCRm0Oz9af
rZl/A288NqiQY0Sy3sfpCClZYinBSsW/sxxde2l+q2YKDx4fgsSIiOxnjcYf4r5OvlSPG7nZOpIU
VtV6DOW9a0ekuuNP6i8RyJ4dXX+PSIAwMABzx5bgysRneTkd+UNNQ0KvJEVuves/aHQkSHEx2Hln
H7BfVu6DwUA4Xw7Lxi2BVkD7CoZCmQRLQN5EsZXVRwXeil4EvDdpOpgxzMG/7e5CY27olcmRk65e
t8eD/gb98an1cZpGMPTNhLTT8KpjpI1esrFa3wC6AtGV4XskgFJIsnzw09un6akdDYxlCXr1VuKc
iNHk+9KfFt2Y3K3HLataOCvmvTHD4cnK7AUEk+s5teFyqACjJTREpOWElHPq445YYAsIZ/GuLrmy
k+7LGe3H+lBTamTJG1l8eH+nATUJYkdCl/teTd/juLC7One5qH/L+qCukWrpN0vyMb6sF3i2rs6q
+uCmEGWdyS5MK+KrOvsI5C+Sy2tbrFoFgLgPzInaO0CXBlhq3hA7tKAM4UPG71tvlpMVa4nk52gA
nMfi6kvmmHOdbR7OKq4k03HlnV+IlXJAGIqKyqZ0G1RWX8PLkHcfV7zJeaNt4mrECYkb6Qlb0ov7
lfYdOxqyGJYf8pMmchxHffYUSTxmvSxuMmEiuYfix1odtJzkdsSDh/WAOVw+zQwzSTO/0fFB3Kub
kmItMAkRGgoRlTp4LpIVpc90G+tK8jKdq0M+aWMbO4ONPYJ/ZgwHbHINaca5ScBLrP+GTax+ZFPb
kxf9IGzAIY7MzXhAVxFTZ6uz36y3v57Fe/nl+77exrCLrELxtM6YRXQZMLvPQG7kcLIYwM89G4WH
YWR31fdyYurIZJfnBENI5A0HiWIk3MBi9VFc3L7oLEXWdmxqBkKAANtgCxGKLugjFUkckVS/Cjbr
IHIa5V+Fnbyn7Aso0bo/t0JUEGjTDZ2bt7q3fzjFqVQjBfGoNxNsU4G6HOs3QDGF3MNOb4SON8z3
yTrJpeDR4De9o2dJNWQytnhuZMWDN2HJFo4ZnEPvdOT5W6vnTEa36Dkdt/yljVicRH7QG4yZNyYR
d6/DMmvdLmHOkFNbKBBJV5l6zffo6qa2F/pqjxCPX5KIredP8xkULKCL4ZH3AfIDuodIODyo4Zcg
xx/iDVHkbW1Lulr9c3OgQXkwcnRPfh+V2zUtA8Ct+0kOJrwInk8TudNhQcoRnR7KU9HUpJ1dO4CF
NHW8a1Xwvaff6lCptnZg97HZ2L/OzOMEK6nHFFtHHMZVNzQH7Ks3F6fFnjMnzc1t6T/jNerwxc+S
71W5PulLvKg4T77bPFOMJmMsgOKS+U6skWVMuM0RA97a08HrtDYwFWjytneARU3Ywgwte75toEqy
uAFwH+fcD1l0P+UfvxNQEvYb9r8fij3pXc9tKLmfFYmPvA9z+7dnoSw9mUzZXwLdj2NNgvx5v309
DO+F8xptDpLkEdTq82GMHRDI9Gdv1gM4WSkFh0EHnY4phf4j7AKToKDXmdWuvy4U1nNn1okYTgi4
5MZXG6tBwHLwB1lyXrjai/7EUmKAG3U5qwfF9Iwxoxdvc4LwmhcqoFfRDuzspmL6hIRXlcjJozNT
HS4nw8NI4DaJHZvX9oPSlt7ul4foWsQpWyiCRayADeCjwFNBk2kryKaKJtQpIXgJ7AyVoBVv5jux
/d4XDaqh/bPHzDqwgsZBrMB/wsilh2ufKathXV6HSgd7GNOrDkSK9ZXffxYZ4TlrIJIaY/HwuH9h
C4qKApfep8jXA3xCowkxWDLG6wHrbDl07RkqC3stsiIOG3OwA7o/d9l0n7pWXlmzzW1l+/So2Fek
4fTuVd5NwjPMwSrvMHCKC+GY9N05MOcxsr25iqHo6Rdq1u4wZKD7CkQa/yVIz4iEfsyyK7TJdwsI
oSNjmwd4elMDRDJDXmapllHP/4WVeyxnfKkpBP5gZvA8RFH7kjcVwzOLbYz0zopefgc8wxzbz+n9
Ie9Yevqeuz7x3qm7oV3qUSKJkqJ87t5+dXIUxOLwSnNwayUYUidAfBpiUswnFonwTXy6f/wzKHeS
Ka58v8AFiXna8S7Bcm87xImHZe5WoxZRiketJhCIwCUyoBrstgSYWhwreeubLGgiCpn/gaVfFgC+
zwm0tCcw/Bi1zxzhAdI1GBF0Vtgx34Q4ZyNMBo1Z/RS02y6c37nhn+4zP7Jt5n8+vmbisPLu57PD
RRxqAsqdPGQJVUayKvCfdGByDi06lJB2NGDtIVkuP0NFw0ii8acBfAMw9eKax/5D9441GcsNm1tK
XRfmnhQKcGgIER0useWejHapyOvKcaNp2tlgKTOW77gjuwRRZ2CtARhLoTyy5ueIzXrt3SrcSXhD
QpZBjFrHLCQAcADWzRJcW8Ml5GBIt8RM3eE4gsgAGoSPvS5N9aOiOnXbjPsSpvSOKSAb4UIKwT33
416U0fZqUAZFE7On6Cf6IC8Dx5p7o8PsIXGQCvZfn9xUUsCR1mO6Mj/7GYkhuU46yMzat6IkHoWx
Dv0JO3A2zArxntMXyp8BHpPBfOxoTGymAC+xmfqj5hk7GscPFQrt1IHSTzf3NLVlRgqM9bpQ75Mx
lEq/VOC4cNY2dgrFOo0qry36WahezqC/Yw1po3QwdqgPPSoSPT+X5/mKegcIpgYtiDjaWRzensRh
tt7JVQKlzHiCp2Zl66xCoU+fQxtJkNTszB8RfREPjZmoi8qHNCE8Z84VOW6BwyFsED/Z8JIZG0/M
1ZK3d9h9makG0A6/ZLKUuqSruNML3EO14SO7H6c0ieZlmxK2odzHhm/f3351PsaSS8x6KS2nuxF2
tmbc40uqQKfMEhZFteqsEtOudiN+4pDa4GHl47KS/X4zqyGKjx3vfmYNStGWe5XTDpyKzLQLAnIY
aBKwsK8k7xh1LYrTsn0x9jkjvTLdSOue5/6EKDJRJC7y+XbxiaYl5yH16W6nCn3cTRO8063Y0fOn
oQ7XwdY8ylweTtFHa+YVBSual8ZVFlxleQjPlSetSwJifTnnSA0qVJGfRzx8UgoTdBv5V9Lip8OF
KA389f37asYONZGIFVlchnanRwL5cE+u2R/kOJJGukXj+wwJ1bUTk1F74dA2U9PwDAqBUGcwJAs1
hm8QCKGXF6ixJteBeQnJBpaKTQQNIkLsudPu/qSgOzhWoOdH3NPIGSDMhf3UPTsk5UkqeZumQTQK
+7TBz1pEJJQ5KKWBZyO3YPmBGL9iIPxdpk4DKyUNdX6uCnrDgmbzTFBMsj1ao/Etgxhs5MrOkdpQ
R7xi6Wu7lsrcrMlDELIJY/vdM/HeyAFB61VpjzkDGdWcpSc5ckSgvJLd8OaJ8hvhPR4k8YkwveBr
2ZGvtxBqdFvjz2q6rDUnHw7UFztfop5t7YPYenrlFuGSI+gSdFs0/s1sGV8ufhrSxlKJBGKLPPVu
go5E6ZRLM1NuxtzT9aEvDkIikE/Arsu3PwmzRkGUMJ/bUis+YDHQa+9a32oRc5Te8l6xcbvg4JYe
r2JRhmb1pPH47ujl8iMVIIct4j8k9qr4cE8aWu8weumayqrh/GnvWkA83rbVOw+VLPbd1WzFqwtr
49lGTzj4glkO9y6HfrlreVElXpQo4OG4mPntFIY7ZD/m6K2TlaLsnUW5qU38WEtXe160+gAIENMY
69Cnx4pUldInmv00YPNJBD8jxL8DRSsYkxAlt0IiA6sNidyyAtZIykcsIxc8LMhbIHCvNDjygLit
ENyuLb4W5kDs1x6HBeiUa3vjNxUYwp7GW8K9CGg37/0inZx4oC7RV21C/q4exJeGnBeUcnZ05hxL
ezGYgvnn8x+usJS208vm4OXIFcFQxVqhWDbnkP6Ro0amjltLMMl8wTRizqHKuP8nt0zG4ySm0oKY
8b+2xcxpp6SbX3WJxSyRXUvd6xjOh+xKwHlLpEa3QRnR4X0NI7aQS3Up0o32Qmbsv+hVp+KYIXcN
PLWeh+1Lb7qGHzXJzot6s4v3kVjCimq0LlhU3hclqAEok0loHoXgoadhuU0cfHHbb/lFk3v9SENe
b2x+WYrqhKo7xkI2hsISPZpUJufdvGt6CYteZpQDNCVz4LXNyIXCOM3d68v+fcRbbpRH/ThDTjaV
eF5z+xnKRE2ct4Kcq3/DNihqb/saAmtlPU6zpIUWr3cBrfxErsaZ1mMFVFpp9WZaWD7pJEcQxoq0
F3OsE2YhS8YUlZQ5wvfYju6J9feerXE3U0yq+P6vZS5OA7H04WmoBde7IyVoGL3meIphYcoRw5BB
C07DSLKChkymiipCde9kY+EzugxxwmInIILo0gzZkswnuDv+HgdR9Cl1QkStCOrQQlQnw43v4vsa
U7723ko+0+/VPxH3jVkFDKrTB1rXlFUPQfSCqra7zfooodngCvBHyjUwZ2fwkhLkO46PryYnYD5+
RDl26RJGJd6XHXv8VcSrIBnA6M3mzQqIXCWYCsWCAkxIUjkgUFJ6+YSA/L+6q334UB1S/4SrR0+u
zVs1ztgktJYCwA/giVlJ/f5Ikd1DnNMSFxn32shvMYG9ujGPrR/B6DsyazUJzt46o14EvZWNERO8
amqKVoHydhOolvNKAF0PwhoQF3WLZtCzo7qpV04oJiuBavmoKJN0yFy4xngM2vdZpN5zONxDHfIJ
rYYTKc43Yyt8ZUyzL6Ipl/4TpJ33f/Kv9oYX0DkJHHKW3lnXVtuKdui58sv3APezL/Tfh91vU8Lh
2Bq4Sm8de8Fw9jZGv7sVJI3dh9hehIQkmvem93pwBHdu70ykTuSMqiY6wsKFt7zTsjcJxWlTWMYf
zRi4o4iIadlfvE3yr4wpvG7+xxfoU7WiSoh49N3mLZ7LAS7W1GDHw9HJBhBeaRAmLvUPfDl2v7A0
t37aWWHWfaYd57J2exhd5XV6JxM5LTu5ck/dx3MV+Gf+3MDMRT/CZgTX3cxuTLaP2JaoplxiBHgw
y/moUBZMLDBKhmKSkp8BnU19yIuFGFL57ldzVGj5jmo4U7vBzCb+G+mom+E4zXVjgQD7bgEGvZH/
UXda4dcqhOXnTb7+bzgCZPsRT6CmXuuvAkFYnLS/3dlNwY0xKZbkdfhw2JitRnzHro1hxlFoqpm1
yGQPmX7K92XuO2qLXtBe1ONryuibnwlGqvmnNAlmzqBxpw+sWW0r4I420hJoLKLkXOvHJykqanb5
/J5Lz7SjQwqPKf/cVHxhT7sv/nFkuKrgCXVhC9M9yiTDDdvekjafmizHOqsQg0+Z2L+Q7SIPWCo3
m57VqqGbtfWkedwsV8C98SajMIaEUzuhwl8xr1cLOc3J4Rl6Rh2du+zw7u/f7pYwCd+e5D7hBysl
8EgUnId1JrtC/1jSOCwzQJtmgs/HGG2IKSepOrZKkHpOUJi97UkbnTh4OYfuIthhgTOFZig3n61K
0w+QZQ4OpVKwDi3ARzNS6I3BOJugxl1rG3Ly7ROzgsDNOr50/2siOUjrOznEelmVrgeEE5My2/zM
fusecqfQp3wfacvk8t3EvxeNW1TxmrSWwgYDQDe68TRJtvjDZF6NC6k9feKWb2alOpm8h8Q7G7oA
Tvz7tvAhR3EcCdav3dc4LjrCjJzolT+J0/Qz63IG1s/5F7TKrgQgAJRiyogLYWxVWDzC8g4OMCI5
j5lwWekXWAouXrTkBZpxd1opGguRS25ITotHbNSl5Lk0GigTLVkAVHmN4a2Pz/lnbcIq1I0iOrZM
TWhA0Z4yUfUvsarY0Ec0LQfzkgg/ubgY7EK+qo+0yEcYYf88QkDCOO94Qjy8PedK0ioyCHDalFwi
KF/z1VVqru21Yef37viX2UGsgzsRkLfJGwcgf8qH7r6nKuu/BFJDxIYoa2Ws69xlhHZfbn9l1DKg
SaYKORvWRKxl7fnP1zlncKmKCCnN8nFctDQmAjpWhp84ips0lXSzWkMc2wRvZ2jQxK1a5LWxRdVG
3ZSqc0xTZ9W3cJXtT2mNC+fs6QLFjGxLaGZyb7t37TmXJNWVntfacKvRRhcT4iwsjoV+ONRN0C/g
ShszG9dtqvGQbbAcXQtzp+8/dCxZotJ66iWm4+igCY4dmzV0sCwDOXp47T+w/6g9fwIwuWP85EmQ
RdfCxVdJZc5dYpPxV/fPW5O/mZlVm6NdMO63uStH5vqOorgNxOv6P1UKJruJeITpXw7Q/feLyKjy
YbaT3XkID5NR2hVP7SbcQelDRvAEQfPFTLLrV4QFlA4GoD+MMw93XhQDBRzQZaLG+Gf+u2Bh7cN2
6WZMXYOwXsjO7xG07RBkmPfBPzIFxb1yDF99NjcoDNJPNH/G5yH795uNxkajek2IMbRUtcdAaTkE
jjdLoNLpCU565ZIL4QOW/ouD8z7asimRN+degMRzzy5y3iiYG0hqva2B3YBpwJMrRNDUeOhkhK7L
/iLNSeO7g/FGJtksfQntKWxskhhz22D9ZgxSWfzxB9/aaqW+BUyjxzh2f+RRzJfuY4yyQpWIPpQ4
rx07xoE6EA0ANJIlWWo4vbXgFaumJDjDGAcZg6QaoIzIUbqzn9sgLRVAS2Xw40iRhlN0o1u8XLyH
99xetjaMRsOtvtooa5o0EOmLV/hQgffgVimCYVnYYycBTP8ib3L4LBe8J9WroTCGnmJvEuD4MELY
zGlFUBcBBM0Xa8DTaIWkI5nvfwSdQv4l/KYRj+hoxL6XmGLP1rePLHDamyyltz6rQroeiM3o0URh
WSWcqGhuOuD0qjUBozWdObkK3EF3pRHl4sujiZ5U4LVz7rlYQXWUCeCmLNaVvDBDOyduKcXcWC0/
fvOEoGpVZzDIfZi6geIF6UczFJIl7yyPAItAWcENRq95aC3H1XOcy4QiuHzkZV8Lf2GoBGqffggN
k0Luwyklc4YYsoAD9pTB3x/skelgfui9qE6rI/nMiVSdgVZ1cV6r4Mb3tZrA1Z+7CTyO7AlZU4Rf
chBxhVqbEiMRDtZHF/062PznkUQ7N4eln+BcgJpw8L9N3t3MSaQzA+n40aB9n2RK4oMB/nAEf8oW
jdCeaD8f+Aghkzi2P+cc60uxFvXBlSeYMtyIATtVddB1DcTNcUDBeNNTl+LYe/q7Z6ZFXKVMZAsG
taYjYbdFAlANfbrmyDSlwBVEbbdQaby8bvb3PoxxH3mNpUofMclmfx3obbHav3a2KrGYR8zBsTDx
K1NnfHizWQGkQKwD6f7sYXoadrxoB/MMlZ4XkG6mhWivDB6QyrThdJ7MmnJ8kAXiui2z0NGiHN7q
NyZPhjhT6tOCFU6yJ/yxHchg0H+hsuzcoIjJ2voqAGIphLi2WIR43rAB0NDfPnODAUHvo2t/wRo1
/w+5106+RU9v8yuf5+bSAnZMmktxpd+BPNktk6PKrFMd148TBixTlTfnxoq/0M0cky4yYQQIcP5r
0C+xUeIVPtIuAjD8a5dLFHMm+yTaOimokhnXTBh3ZnsWPf73C3YWlhy0FD0c91dncRfUteJfXe/k
QykA3qoUVus0glNH19zuuohuBkKiH9wj21CIZZROPg6RnFx1K3z7q7Rebh1md8NemZUJ44MTq+Oe
dIl3MZbdDaNY63GOEBTH42Eb0+rAxgJVOOic6j5VJtb5LvV733u2YpCT+N07Lf8p5M1D/mRq6bua
gpkCchVZU0pe1kzIUeWsXZ4obxD2N8Fy9ie8kS0t8o/P59036CbfPWlESiEZrJ2HgxRSOwf2JMcK
e7FmqBP0bEW44DnVEuygkjvhRGNBUPZyvm8MivcLf9crr2yPKAZ2613tj9sQgN3Rj/XCbwsZn5j8
INxrTMw6qt4S0Zk6ocSD+csAqZxjJz49Kxuo2dAWxZWkQjnUzklYlz8RwC/Cu9pcmUVOLPbkCb1d
45JpURqdE+Z5l+bOSDc/XEg8ys7Kx3Gl8sGBS1EPFG0HCkOgZRTtOuYA8OWbRe4CW9BHH88eefu4
ntegZKmj4zTONyyzV63qtFbJDYNb5HfhuBfE0jAzWUp9Mm42e0e7ML1vtsd47W8VTL0TrooX3/LC
1eA8zuLROUTUXxHqIHx08Ug0l734DV4lvUztZmGm+xLuNp/c0jiWzvyEjGGhToXmOCOES2USbtNK
NzTYCkVlWj6lrfb+qmF1kflfFNqwfIYAgbCS0e0K5W1V3JwtdbMKE4ypZY/RsoV3ac3NOKt08pcL
Kx3HgQZ8to+d+F/FIWt8d5xvA8LPIZupTnbfSLjSdRa9kJiHj2cokNcdinVQkv3mZ4aSFAR/eVVV
xvHaDJMbvUwRdWORPrJusDnbe8W1UgH5zotNwcs0/gu9QhVoNXaFheJ2iNvvIcoxTAM3MzPeq1Kx
2vVV86xjpHZwTSvXBt61kfRKaRe9Z/VOw9gouJwfYPnb/Chgqaz5YdyPWvDXdY87o6tjWyULRWi3
/MrFlorUFJKQFXXSKLQ0Fe0sammKV11zM75wdiEhWFUrwpJiauVWc2D1Yj0f24wrsJzkMiow8CBU
zXPvvViq6Zgr1U0cxsAOCtOpIqQyQYY6L9GuSP4JY0WbwHYZouAUDW2m+yNv9JwrKmyxi42DFAjT
YEq4MiES7excrIncfxhLxnX1xoyDGECxw+mB4YPZBgCo6ee/teLVG9R/wUVmTx9wl0vczRHj1V9g
sLuqU3YMrfcsV9MBDWRQBsqVByfTRdc2OhWx+Kat3X0KoA1xC6wQylHki+ntGjgnPUB/t0P1T9v7
knUyV/EFlw9wBQrqYirCXAe49PcuNai3KufwUD2zKH242L1mwJAcqp+hdkLasVMnUOTVc9tit9xy
H7Dx+j/kkZjVKGRCw++CJeodCXbiiyvGZKM/krh2NirRSn05s6y7Z40JzWqoHZC2tDSyZOsybIbj
6KnA+s4MrYlCZl8yYTbQ37Z1TRJjcQs5zZ9fNCJ2zAtCi5peaH4Bt+Vh0Eaxg/LUv1CugEn2v5Mw
mS5tTVky/BrkIBrcRA2QgxVHvqB3YPpWMHGVElTtp+zY3T1NqfyD7NcOpJIFXgkSV6d7zeOR/VXo
MU8H7LT8zOfpdek2v9/uP+0gdYc7QrfBtw4t3aSW96N25EbJ4xziR4jzQ5CCPzaEP16ngeFkGail
90CeQ9gMUnvPdu/x9uGwfevyobiv5NxFAuby5vrvJqXUckc9nOSQvCJxiwf4DHFizt7jBpLCauz/
bJtaSa4BrNic6rZNA3HeSSgub6RVTakrfdYojkY8gk3NCx3u6/TOTZo+WTaySsU1+w9qHxwXYzyH
kTjEXpkg+K5Wp7KHRNF/YdGiAkqKkvyzqhyRQuM2jnefNxdJH0lg6JCOlslDI2aQ4QeV1W0v7Tfz
kJ+JXeiUV9dYShD33tcr8RcdUjoO9BTwFwPZm+5yfaR0Zbaa0VCukJQ+7S7biD7Cx3pdaMvzHjpC
iRqiryZ9rKFoFLZRX1zEvPtygWrmwy6/e8nfXriB+jzH/BecTwtBfhQZfNjrGRS5MCbCxcqtrS7q
VJrYKkN4R+64yy/mw7rPyl7U9RCePvXLM//sQIxngGhggN6mRy22kfyF74dxPgZaZDGVa6dFnn0s
mEZ6Y+BHaJNYn8pivydGkoMB85gPVJojvmMPlQ6gXf+nmeNjB7eTzG7dlgvuS6ZHlNh1DAEvF+4P
32QapLSN+qz8DihkIBypQDScbPBrnSt5gKX5iS5WhTmRJ0TNeoDYGwtbGFpEckyQvVuqtv02BKTl
Pjz06STM+lJbS4P425UWydnZi5msE2B6KhOimF6NGBTuMFFh0aiZSmgilYIfqJf3EOTsfStXDTJ0
7gIEDCNCQtSUos4VioH/oKjiFEn1XpsqYd7JLF+rlAP9c7JbS4iFn3i1/dhutTPz2CgYm2rFEn6t
Snzt1ClGpwNHiUIIV/XF+jIRXrydCXceX/I4NEHtcw/7NJAWYNXoKpxp/yc/hmhBhZEOo+mTvS5+
wKdD7Fvmyr9/MdCZ23/WmaOzyFo57+Fn5aVzPAjlL2YxB2ofobP7f5QJbFd0gUhRx4qrGlBIo0Mj
pzYO1gl42mxkrzujXOAB8QiVdv3kwHl8KYhqvyag+Cdf3SdMKRlRYsIuiUu4N3l7EpPr3Ao0ql6i
XAHxTYGxQZeYuA0NnwDMgKIYgW0B6vkLHrWJy/obMyc/gKyna2+4bCgdqpiLJqiBQU0l21IkuMv0
qOu5wkYTfL/olXfW+W1U86EuYXRNrGvSbHYEaMDHHgVzAPzhGNn3TCXDQniRiSKEfJ5DS7ERzNMH
MgxyfDH4lDwH5qPNbtMHI1vHAZ43Yp3Sd5kbhZF31Aw8TfF45HDA3LFoSl8LR58k7XSGT2VruHxQ
6ptLjpKOj06r2XBQz8N9kbTxqgDqwqCsoJOzO2uTnkRhvOyII9gJdeyc4o7E5SZL1VGD/qZYMXyf
5Duni28A9Yy9IY6u51VHZTRkS/8HNaOVrB5Mt1pKfppI7XfbHTe5loQzgQVFCROCFXAWJXSslxGn
X0JyM/QNymovUy2W2oeylnXlwQTa6u//JYh5dI9p/vS0XBGUttHK1xCWxlcarGIQYLVblqso2c5C
lrJAIH2JRCuH8ClT4J+Z3c7NyYIKghy3wOSWjB6ktntvM6WFLvFijl83y153etQHKSIg3PosFhSz
qmJq1tzJE+v46AN8+Etnf8tDx3Mdp7Ha3DpdcT77E5Vc+TDaVGsBF9UtJRP7K7glRDWPY+ps4QlI
WaQIZVGGaunNU4WE2av+Tct+rnBdiF5cfMq6nbdD1RebnzQXUjB9qlvo2AoRnqjLFe3dl2ylMxnU
o8erdS+qt3uN6Lr6F0pIa6eZzksJMuud318VcfBk5d7KvokJ9O5bAo2vqVtZVdxwTjmrYGKlA5zc
/JMXJyxpQJjDIUag5/WDjas8VuWUtqv8jXCtnzT9PjQpodMhAUIrUNjll+OftLxbIz2HrnBCg1ZC
ioynN6Uwrz5bKgiTcw2a5ZgEvInvIoDdefutfreX7uOrNrjIYP7ut/sbYUWAUY0aUY3v8LIIB5oU
SToFmwmaPq90chkdAM236od0exnyvZ2/Z4er+zi5eQdFFryQ3IFXPcSkz6pccPFVQSuGhekIivRX
GgF4WtcU15weKZil9ciwtJnY20kItHDSbdVgVSvOgQ6I4j9fEaShrLhGEWR2jBHvJ3DAHQK2ufSd
OLAwiQCwQrAeSXUf+3ca34E7pCjhXi+gcLvzOZwOnnyvTlrRFbNdf3JtGghgEwK5Cm8P5L9yr0Rb
muVYPxY7xssoe0f7StSGw0d+v3hGMdJItmljQQZATldUB52qcVsBAiix2SRhBTuZtl7/LYjQMRKP
ci1be4KDAG+5fzYPnb6bPyLOLAMFJW36Yd51ZI8PzYnV28FM38d20RiTGvnqy2OGLWhusbBDNlfL
CpVFFpb0x9n/sY3LyJFt5NQoN6t8gRz1TVLJGOcIVZF9cQqUEkxkP0tFOAoycvT3wBIEuhkn78eU
TikBsJOKSbc9vpD3fZTSI3M8/spZw2T5gmcsBp+7fgvyiFNdVHDsy9BjuRZkVoDaV/yuzaAYGqHm
9QXALDH6K3gbppuXYAh2DSXtUl3lDUcDPHuAMXMGLeCT4f53DBuDVSl3ZrTl0X2sA0fqP7TYtBnb
sO+oXUsSS1ERJxxolnGykTaNv60or4d7GQiWOWDU2Z2t44h5G3OC++44yKn+wIpSRkH8OUZftMYQ
eii5PYf7RbQgG4RdA2jukXTwY1nwat2cWpSjl8tjFkHIqeVm4PFz4Nahkr6bo5jFqKdQn6gjVtWA
q75TONNoqrXhZQi9YRbsSAVgdxrIGOtEcWqI3Aqmp/Dt1yHMKvZG54XgKeCR39JVY4Vbpjuw5YXF
sHS0LTX1LUp1bFv88d6BN7bq6wkIpPruN/H6PE7FR2HS0uXSQi4UEkFnr1hELfzJbk4QMXeitxQD
RqNrB+xAg+acVxfk0Lb5EFG1Nozt76Bq8vUs8I8PqzvD4HrFPns9uEgEnXfwO5kY4Or+DueKHyyd
GxNwHAwq4/6SKZLFvrP/sDcKo9vPJbngYsQqSOvux8HJuMOeXyIdPwmbxIp3NSRClKW5XVdPKRmK
TjKvRl0EmnxTePt3+1R9KajT8pRSoXSZwX/AhoxUVdfLchTaYmcIBaycer2WlHEXBkxzL01mnqNa
L7uH4PhecnIBEu7tJ3lsx11Q2YBEEX7V/Y1q4NdM/EQjnyxP7xx4GG1XNhiOhWg2rhP8r8swsBB+
mUFEjW2r0nknT4W4M48MMYDJcl8x2CnF096lXJILK3JAO4635/zgKarh4WHzGcailODfBxLlp3WK
juYqsFbodgf6Lx4X8pDDgmcsCXrtM7siXDduugOruWTdaeGvHlQYwfcR2oxZHDV/d1lrm1PbQyUX
/5yf9+tgazdWCUYrCN5DbpOBTS/3FsXeRntAEyxbJd3/QHI3zW67ARv5W47XE6A62pAnhxOJ3QUK
Yfyx2Bf/HCL+9qdJdsL/YwN1RW9I6w8J0DaWHxJ0UWmndGmLWPY5soY3z/BGKCzziad8e6BPSkqA
UK8GkckA/TSAwLqo/XOp3oNyc0CU0b97m1MH5qoWryAiVPQrZFMgNcoYqO13eOXl14V2X8PhYG4A
oMi65wHUiGGm2wWjEtPIBhy5K6QGfkggQjCc5t7QupPA+SlWhp8xu8jaD1qJri/4iPG3Tl2qIXVL
2Gt0sS6cC7dMfDLGkhcpUOsAlLkPN5WVDlMOrxgMVVA09z9q4HRcdUvWS2rUZs83n9Ojc/jinHV/
2p94fXqcMQGeZC6Rp+Gj5ySPBqWXMlzq8UbxE6fdYcTMDrJtfrotdEwCj9Om5o8zylogEmPcp1hF
zEBMZCaISToQCcqWF6jQmQM6fQMNgR/SwOzkStEUh3553mvtYOIfJJO30x6ufLZNESz5X7DXrcLF
+z1X/8UD53+KRMQcaWKmEGDHZmYzOvtbxtDLaWmLlS6ZxsRsAHzO81ahJgfwjgGKKrSSquZQ+Cjz
FVMqAvTT4HY4TJxBRdo26+k/AEJM0fztk5PbddXrkTid4MX90y1u7g+ZMcgZVj2yJkpyS9LmyoNF
LG+YvlJCYywr8g/J4gnpkZtDT+3E2d2xpKeGdXYQEueQU9qwheGMTUqkLPoW85ul9nR4nZng90Bz
fwpPpGnQMdQGvoqXaylXbwyrKTSdU4oGiuxsghHAbfFCDLbL00lmuXh9PSWtTWH5GmkJ7nC+aKpd
Oxf4R43CjuQfbkNo4C57teNz1/MoJs9Z8sp5lW7zfWdLdMzxRIjM03DK40OGSezq1KufoBjfXm09
UMfXu8rYMCUtAbBnvCet/SSjQnMR2oLcHv9QXjnElTrOtqP4QIc8B6gkPM5ZqNnZ6IhFi7PyLXB2
zJhOkyb/dWkdJCiPJCLvIZquD/RlgTXngbjep4QuTSBnNtKgT1WUDYCXU8Ad25HF1Suoy6V0Ltor
d5sIDjHICF27b5SC/r+zVTNjqsJsUcMlCnaYrqFOYEJvpbqW23EVrysFVneu2cZFZgtitvWttUTm
1M7FsnqNKombTEd2EZj5a0vc+B3eG41qz5s3zodxK/AcWUMW/sedO1g9EENRPY0i/AgOMLNsaDhK
JIf/81gC7Lhwrocs2SPBWvEE/nxMkAj4+IR1z9hkIJ6qm7O0JU9VARA32ireKWPyiwaV5OTZwnb9
mqXldO18gPYCrcRM8/3djRd4bNns+FCMnfoy6GNT53kBqv1l9u8As1pyfZHQv7O9EnE/H61CvUbt
5JxyDNhcbkf84r4YqGMFVEU1OYhwLpu/H2HyTHBXwHopNP80/qp79DngEYE+LH3tj1Tzo1icqKUr
XadtZcHSk3+Ruk1vTU+M86JFfJLc3YoLjwRdqJGlFidUg8bOmy9Ytsrxta4DTSnS44V9R+Gd9LLe
VQl5qu/2vCdbSgeO5xP2CzLncRDZvSES5maMsGd8tMtE5joI9MKbTuimonzCtN2bO/eelDDMk6S1
gjHZC+HLbqG2jrdHWgChc4FhzagHXpAiKs//QK6QoRXu9994jHjCwvtyAqGIP7FYkyh4YviOxJVk
kN3CgeEic4iCqUMvfiHTzLrdHo9etEKwlmUn3oUuA4aNjWMQeGHAt25YFHb7opg8Th/b4jYOKjg5
2NcDQKQGPS6wuSQP4OyZZdr23u+zOz5Dy8DsssEw/P04vE9AcmHafbDjAyLCru8993cBAecjOqGu
eoJoOfFLWOnDfcy0NDuqLqK8/dSBr8OpQUg5kDSePrI4KEl8zg/jSSlCpqVgCKIKFn5aqTtW3bao
5/AyPl2j2dWzDJIuyzmqOgJxVdK32eDfQpwtMPVQ2jdEpXbB8iQNOdJXvJ3vPqdxAYwLXZ4xMs62
wlXHG50jCrpAp1rPS5ACK1lmVw3EoLfQ5bBTbk1rDciYckAsdagaSFwQ1ND2ci/tWqdmGvMq0e4M
zXYqMOKC0ZpKJNCsK1GAzIFUN03HYo9iyj4BGCMYg9xg+BU6X28NmnBOR7mLxgRSuJPHlH7yXlNs
tvPYOV147SS/tSryksb2jRJK9+7jjjK4PhYIbw0diEx65RlN4saSQFilN8z2KaTEgNcjWfCiB2bB
8JsBKgV5Zg25ookL5KY+o7ez6Ns0YoJp0nfVEe0cba5oaYnhUdK5x0jWH7pc29W4MBjjrN80sj0j
6ysluwdz/3qH5NUtyV9b1hkh41hBVp+aba8r+WyEgFXEupxHUuLPSVDOU1uJPgakTCXCHMQWGr/y
7bqPn2OMcFSwYYqG9us0a3W0a0+98Xc4hbAfF+eFu8CmgXj/Knu6fSkQlqhMydtj4t1K7lOnNbko
KleeoTa3j6Qb/EO5h09vsDkp+LR+HIpFPL9v6d/ov+/8tRbir8Tu5L++p/Sd57kkjCVgFInAm77k
9vOV3pkSaNlEJ7u432n2IPnZ0wnY5wYRTrPnnATcXP1nZtjn93Qq9SgIIaJxUGvikFQuatmbzIl5
GncAaYq5MeGdWZMBNbCOe8zhAwGlS0Qldkce+wdzbGsfjF1nioWlS1ZOGkGy8LvkchmHpM/Tx6Cv
esh35oTJ1fr94iiYxhWyc3LwwSif6QEqe3TeLc14Jvft+PpVr5uWHueNaA4MicUzlk2/diBiiUMh
s27AmAaiAnaGyhQgz7BUxwDIZf2/GBWgbEKgudgjQT+6YuBeMp86UOCXafFTU5qwRtoM2+8y0dhZ
mqweaht9kvlfuAE3P0SLf26GXqWoEvJdpsb9tkhrs5CoYqoQditcj40xzfHUiQ/43MYW6c5npxm0
LwKowV0N47dkPq2Rk1pHkg/x4UQdiEI5kKh082jI/9OMIkHhFPprHvU5AX3daT6L4qz0OkEj+2in
EMdEEXRZJxiyfeuhjuLcB5S3/sWpX03IIanYBQIpO+RO/LiZoHwh4CX1oRsH91H2PU9xm4OwufTt
QIqeF4WlITFPSoeitkYpdlWvdzXtBTZ1yj/olhIoOWFx7qzj8TtgoEZbnh4AAH2CGgvA9Bgld0Xf
fTXIGJdpNIeHSjQ8L6NEJQD41uKY8PadnpX9oaPcB1th4rEImc0Ax207tmm6N/BJzkNns3UYKCkw
GbLEIRRynhMoIZE57hC5hleN6vhtGf64++uvTGNgajSx1mach4tJn1al4d8fVH9O8a7x2go5ad3h
XXW7bECKfZ4FE6I0aDL8tAp2t/kzTGMZgjeeWDsY14hMGkumgwHaxvLnMQuLJIe0sze8rMCxP4oD
XrUecFhkPpKN7NY3ercplLOnSZzn6eiCmD6EGgK0HR7Vp9gJBZjlcDb4KSuhX4I/zUbJM0GDsjJp
Kk58geMxQ0Ucfki/Oa+Dj4fS99d2VsdY8UvR/goRF6ENwrUvtTyYxgwvxDL4qhE/9d8TUT4w7ZEv
0bPcjtid80HdCM/xZLJ0tFS8x5+HQ4p1bVR6z01SNWK3WUL7BAZM5O7ym4l6s0bXs1SwnrgyQjBi
NDgcH2r9slpqnaJlHjb+/Kmx9xmgJ2fnnspvlJed1raIgCQy6GOkG8g45N4r1KfNnXjnFcuQHFDN
ca/Blzq5IvXyVgSMrx6RY2DGyXKeUUjzn3X2FXN6pf4/HFN6g306t6eAMBYZ1KtUuRo0lMEvmZqT
KkiiL7BZ0cq6bXoxr8xMOdSc/BET8Ud01/evqNgP4fx4vBTUo0Aph44IidXG3Bdd0hpp6SsEE/XQ
7DSzBJ0g0/J+SjIeA6QJdsUTbsEIx3uBZBY+AuJSPy3RRx9x8+qyqWP9jfGxiK628QgRnOTpv9IA
cV+5ynu39OMxiNEvnJMRC4QytANtZGv1saWh2hQMMxuvpiY65pbqfPlXmOVqf9bkVexaqnB1JtcZ
UhYNAep3Tj+wZN8hLNwPd/FkYrxvPW/5VifC9jmqrSm4JgUB1iVLIVD/rg7IiFHoMGFB427MhxK0
+lS/aWH+oVPNl0I6ToMoh3I08p51KiEi01GPzdETdGGYfqCiSOCmBhGkGmuN75EA+sSonrF9D0eN
8QfBNM/CrnRLNs/xmRIG3VBdKGUfmG5hBAtJoY1Y3S4uf9C6u2tkcMVMeHhS4ex6IO2FLXBoI7GP
Q1ypZIiF1jrUaZtm1hjtVAWJ8LvlUBHgM1sy6uEfqReHxT10z88NZSLAG5va3qH2+XuFgvZIwTRW
3hptnEeDu4JAdWpTxld69c/ZQgeyxSCr5q9VS3tVngZ+9EiaMcZpV5gP4Pc7FdSRgDuBBuqcS5+y
PkWXVZEY3ROXGHSGI2wu5/Jg+7AdhE+0wVWw1hEq+mvYKgNCNgahFsVE9wp/j5FkvQ+AkdJc7/Ss
GIHCydpxj4/B1iT4D8DuRSmxw1NV+QmlzWMF4nduT2abvYaZk2Vtuzsm8u5jhJFVvT5XpTdPEyen
TdKQ/uWb/QwJcbDvaQu/hPRBhGc0hKi88oE9uShA6GK7UXZoaoqqthaJrbf3Hp33W/gIKREHJo2p
o5rnpOfsyxqgOAoMkHLUhj1wdZCjXFFMVORPqljdam21LFCGm7bnFC6+zRo7uqhLJbCob+fv9QDl
Kf2h+UfHP7vltob8WBaBUhQoXHKJeeql4oAr3iG+ybSLB/x1nbeMHKhijN/tlwe9gm5lf+UTAeVt
MdM+/csGuCF+zkLVy3oN1IK7pBawow6dsyntV/8z1tffi1s/XapDQlFAEohCZYFzrjkPGuhRV2dC
2cN7TMvJ2Gxtz3sr9GKhiepWOlBm55Lp6qhiuNkO+JC2KroY4tbuq0BY1yObhN/h9wjQXel1bX7s
nxYe2UCZAZxg1nlGW1YeDOxdKUhtUsSoBMTgDV3W/JKfmNh5InFMyJM2HYcnVK7us9Trhfo7abAX
8gg8eYpi6bqatLejV74G2qbtr8+RH7a2txWQEP5+HGhCVcsH0AlAW65QyU0ix5DVvIWWazvoAcJ0
p1EzVQ1gn3m4vTwT8smfYAaGoNAMICNmUPD4ahqiIgLdH51bJ1AqUGiryOlg+/i1/gplwOVQJK0B
TppwxVpolYJ3XO+DSGmRorcd3ap5br1ajaLIyIMrNwdS9yhUXxGKD/TORrwE04T5frwPntfV0V6y
8HbjWSuGTQDI5g5N7+GRVCALb1J29eKJy63dipqF6Yr8upqRD+UsD5c4T4zRrdn0IqVJmBu6hhC9
gyjsHCx2MS650oqgQP1/FE+aIQmvWHETKwzlmZc/w2Ka0TM1DBdbRuVkkVGllYiUiHXx0BxtJg03
Yc3tTVl28WMX50T7WdQetEDGwAS0EXUmTZLNvkyOyAXgWShS1b/vTyOItFacK6OCvJwIwUlqCjig
pDDTx/eC4sw2yLEX9s70Vq9z8v8l0KwzNfn4QtfoZrysSozz0CmcsQkrEp0RXfFg/dUsiTbsIl2K
TT6GydoFi+uP2pj3PAZ68DO9SOyIeL+uoAaN+G16vMZS3sLzFVd7121thXWZ6Pmlu4sT7DpDhaw1
imCkp4p7fb1W0wePOigv4VA0HqQhqUXIZpYaA7LCoB7PIbXVXPCrtue2ksHN5EJzqgonw8ILk1gt
5+GNmFmEmO01/r/To9zbZf9A4DiXwQjIDOgdqegvjpsGwiadEnHTekzWhhQmcf4meH1DKlgmXicH
eX3hywwEZdxM37Gx75sIT5SkwALge1HHqB0UxPJUtC9Vd5tXlURf69GC/33bTVAJpLW2w+dv/Jh/
GMFRTTuwiqmNF5i4mgRdzQIhWRyC9FnpK6oVDTwWRQFydO0DVW0CkpRkkTfRgl6MoadecUgHBlRx
GvDGX2PvgNEQHSbHoqlgvejPiLOUaGA60C6ePuq0uq2PQ/vKz67z3kOBAGMYkrFLSPrYqdy67l6Q
YlWO7VahWTEtZ8pci3wk8MPounZlD8mzoqdIaGq91XEfqZ8WhlZ55X32wWKlUFN/FHf+J0YJgXzs
WnXBxWqSJwJHs2VvVxsAfXF8EkDQgo/7WeRwvtjKCrsQLKHAysCYCgS6A+PIoNWApureooOeO/Ev
hAZ8Ofp2Figy2juomJDVlWK+Wx2VxI4xgLKqzs70b7PawD7h3ZMutMVxxbznCQVI8OZLV/JMHWJD
99BTmfA+asc8wPKLEJo2UQ4nXPgEgSk/l8I3vwU9UonUFS17NtodaC5GV7jCqv8LkbmJOzARgbLX
NExsHfYgAfyHuwNid2Wy9X/nY/J1I8OMTK+hbow6L8jlubsFRbx9IIvU1yuOsbobmUQ9E3O7rBVs
xy0Juru8U3KLXh8/EOvuxQ2yYsXjrRbFHzIYeiXSyE+7kK7/2Hni8kwEpMYSdCyE1R1uApuUY4U7
E86dc+7AsTH9hgPrDJS3IUycdNFhdUkmgduSgneFhKs2y+Y8nFqfXCrurNWcvWMGhUsCIO1aSyPq
/ffzU8FBaRSwhqJxd3b8IMsbR+guSMQViqHZmGepWRtziAtwt24UPz2anfH1KGcFwr6S9ajSRsn3
knuDELkRaT1/MJO7bfz9/3VcRZ9WYtZCrD9vKr/rLRfjOFP/Uc9F8wEjCRtIYOT0bSCZ6WTCfWj1
YxD6yUi5vTCWU6p9E9MM2t+ISFNT2ugxzpC3TqBymestksAdlcN7TUNpuBysBjJr3L7ydsDM7IHK
U5j/DxAZ0zEGhSa8P8H06xfYlp1i5K+i/mwoEwZewdLq+MlzpkuIuzlKWBCPDtoRA46RlTjIvFzS
uvDZc+UbH4UrxaXkqxVZsCOanoD5aeNLitsWB/YZZsiVrTMGQXIQLMweAFZUacfC+lVXpRe2B4PO
MTS3vpW91GRIz7Meger2FyaDI31gxcsrva8rt75prsJXyV9wXhyelCVC7DLkLut/yXcQGDYGv2W1
eyTkFQfjmTL3j8uLQmb/JWi0v2fagjvo9dC6/y9KCt/g4Ui4KlG1ORu/fjuCu7I4Kl71VgE11fLi
rZECDuT763C4o/+r9xNN5KhfQpSqegA3Xd+EkTsuF8eF1H/rluX4T+iAYxXHmwGrn+L1KiSkCaaC
RXSwrHRLckz8cl3dqc5kJsTTajviLr4m0MLg+v0QbGov5Wq9zu1THRnyNEK86zqgSFkcX+4OwFrq
5zrVA83568VxxbO0yqBdvwzplPLFbsq3GGCh96OAAPn76voXYIwr77s/5Qx0QWsWHO9yDIE+/Ein
lmWywk/dnL5vr9a+kICnzaDqHJfA79B8Te4ycyC+trtiTvHo1L6/1gXcVzN6CYDHdOJNiuiRGuiu
QMNeruZUIRY6uBrsc1CH/Yp8zIbzjsWdD6EdfIpA5eKjYS/9/3JuyaLaBn10MZNDiJ0CPTu93nVJ
cawwkuA9SsKnShG/TlL24lTRYdAKkcjz760858Nl5TNVdAOXGTKBL7DQi1O/c3YF0lNsqsHUNMx6
XRQDhR9tNWH8+K0Fa1ZHJrDGhhGiR3OC2+xxNhAbijcVNxROFpu/uHPmm4pVTsUBDpYv/eFOylcA
5WNGLhBqPrgDSwPSFBdblgoUfYG5L/acOLb/z21vNrgnqZfNRbXXM6jonreXos0CKL2duLqgOdaN
6uzg24pmL7GmPqtWrObtxPupgNHBjhzq9kpKycUgYRVCf25eeZjPeFdJPXQMSowshmjK3q5ZWSmD
KT4TD99EDoj//mBdzlYZtxNkC4jxjIagHAd5QrrhsnSnqc2MsyNrOIh4D+fs82jUGxcdu/aj8UMX
PdJMFpbkk0WykHm9hpgPpxPIvlvFeOEWtS4eQGEAXgyt02qzDqtJYKFkj6305+JurHI0gwidvUjZ
fAYDpbpU0yzI2a/aBHvNh+XZWKDdtn1t5BBnFbsw68jV8zBiWFPbfw74UV/MQ4Ub3PfNHP5wjwXe
xjP+UIoOsun7RhE1FCcbJRJKxLtS7tFiKR/A32/W8zUYZTlOWE/OSEPgCWu4FZTkOaB3zh2bkq6A
5y+YojFeM830i1x377T173HLP85JKyQQZUPLplHKGMFl/QqvLzlW4GeqdVWtOCcv+MqyNlArS52J
phTslX7jLyHoomYGq4esK6s/NktuT2oZSFUAgE0V3DIanMdLQnAYHFP8KZA7AVIVPAM6RiDxvP4b
/zX0ac2HwLs16MAWtxEdy8ZP251+C7JoLyPKAHG5KVj1+SrxIAk92XKArK3pMsJakON4ZIx+VxRE
ElYfp/w+3taxkSJD936zCQyK42X+N18b0eanUl+v2sBcB3VSD7KGjrpZFvrmRWvOr5/kab9vQ5Xe
MVqX/Y9hN6aPpJf6DrJ5fABm+dZF6EVMOoDfPU8lKRjdXsnWehw4dL70Kt+hHxYJpyR/478WH2XQ
L8/EJmekz0nWSz8CswsugujrFhhjbGeiOnKOQ+RxReSwkui9VFkj/xhf8nwXFaga21j3FpWUZezt
REuSe2bJcmy3t+1PrwBYkM2JVTuBELkRuegw1bNeKpCIPOt4dKF5UqNenGoU5Oiuy76NY+HMr6MY
Xyn4r6/e2k6MOW+94EGOE/9hJBWxzG5jWp93B6cPIqJbs5yD0SRI/j/g4RfRyG9ZVn5RJ4KMLok2
meO2N+IN7J0iEvFMUFuyKci9jF6tu8MG18bvprXt8gzkWS3+u0AUdqu0Dclhs5R0dRCl2LujwIie
qTi/j/NAhgHXtxV4I1D8zJXPr3VHnRyttAwSieb4vcrMb0hqZ7TMMLi59PvBbnvswRpNDREo0AJl
kRj+CXiI7sDK+3GQyj9hivW6WOAjKMPcGP8uQLY4Dygbsdg+oD12PqaC6h+lMy8sohgJ7pyXXgCD
wz0EzlGJcxaRdZOclRhNakxf1XKdxtPahEnXvdKUTxuPBK79n7qvZ5OqVuoC/aFd+tJplwV2f47j
UTddsOXng1c2IDzCe9LZ+1D6BExCUfq/1p+FVcd3xHxpLs6/UwVJaemMZXzAhv08iCXdfTnYujDT
amY4vykh+xdVdqoG8b+H1NbtsFEHLFfipjzhpFk/ZWhacqi+gnZtqHWzgwUcPNUYm/stwGlwsEzn
LV1Iy38mrtOMetB+wqb0jVxp9lsD6F5ijgmX8aABwQoaljaOJfHHlM1hJO+mOzAuniIEbsZBbtaC
VbpbpO5TwFMyYx8xJavNePZ3AMu9ph77slOVnFpnBEYsNedRgk3+HNZ6wH/zLDF5czktiQsQ29eI
ga9QqkDQXTEeYchWkE8o3islFNREV5lT15qpN7eugKMSuxnGSOP+3QWV2FgXxZNBF4WvDTdZ2Fny
wrg7WgLeK8sKakwjlThn1TTf2qaRnbHT16PMQxmqAXPmrf97l3m7ffFl6uxLtX0eOT+oTXQ+NWpL
GKKffjTG+6nQboIKg6eP3fxiE5pgtAubTixJMYI+xkrQbVYFr7mQsNr1q7MTcEQySypmp6MGtl5E
vM+P/LS13rCSRQc2rcPm/Lig32DYmJTkWnR+PCM0KQmxv45z59amb06I6N1bWRGJI1WAw3E1wOUA
wJY9kI7LbprXsKYgzzwQLVf4d4HBckehAwiqlAHNQ3WYeLc1/wQTSSrUr/9dHAGmCucmBoo/iA1x
J8ivYTZg4NmxWm07B4szyyEb13yaokTmAo340bQUIjB8RmhGKYZuUHNvWJyud4QVmr7iA8UNMLRK
o5PJpz9BYv8dS90N25ZdTpMRlRySJo/crXR7vVG27eZEXkLR+MIf3a92MeVKT+52xvSYCJ0VqsAK
rGXrJ8DA4H6Xbgw/J04xaDi1BCHIrY1wG1MuEelccjl77jVb88hhcnHtsgXtuW8S/7lV+Iwuoi1w
bMn2NkVmMgy5llcg418QIWfc0/4M7nY9L40n6NxCfw8tR4jXm4xK1l0CEUlr/nbVqrfjWF6facmV
uK1rIHIItSLRu6TZzOdn4ZMSdU2riwMeURllTcMy8HAO6tKMdxw1iEq34E3YKgzoEp794e+rZHrH
802a+5/LPLJRmN7BlkY1MAts36e2I7nsYMM1JwBLGC7j5gCWBFzeOGxKJ8TjX55l1vaEy5HTBwaQ
4QfKWotw0TjDMw1oqM2HoQI7bYOHCCgnuOpkvjM07oHrvqR6R8PNRlaYraMO15at7vPNisPeo1Ra
XBYyANTeyhqy3Kmx9mcZcQkUen95dVNRCku2pZpl1Sm4Iel3aK3g5F6I6xDdj8FMThWfTEccchpS
CCbH9vxXyNXB5YI902mWxgrWBEnLSLx2aK+NzKBxhNpKImzZl0XjcbFNsLI+Wvy/Don0YktIGr/x
78KGWI257m+H6Upqk7t7iF8asNjD8h8R33ZQpBsi/fnyC/rHCyGw6kyVFXeUcO/0R/Hh+t0YFoTM
S9zhO/INcudS0fTchyYgkKX8PWr2dMuWVE6uUYsLgvU58QLnYOrUj3lbXhIgDSnswPWU72DkyucO
q7YeIyNxkQK3WIfPhl5jkwdtP/S+J0nemgVElQR0D8AByjnzQIj9Mv/vklTRqvcJr9O/Iw6iRWUD
Sgtkv7CO6OuXPqs2iNK05EI31eFKg7R67psySWj7R855BOq98E/66uA9XGSyOi8CJuTn5K4z89EL
D6IPkWQB9i7XYS5I9xMcM8fHqXsTgQeQO2Y7Baa7EJW4oqo+upD4mMaRN63EWAMsMggUTkL54q7A
KArmzqM0I8gD0ZwT8dwDzJVkX/5+TzO3wAyGgqTR3l6qQKWYf/Qw0Tk3b1ukMWn0PqQAOv2zBNfH
SYZXa1Ah1rL0LASKbz4+tnKoKe2OtFqhXVKtVrb1diOiiklAvDSNOghPGds+2VclBw5H/d56iNc0
LSRn87P+uG+3Sw/JiInrW6Qyu9VIEIKNwLOSnFMjNh3Gb8GlR7EEuI38v2h7JI8jYhXItdAFGPXx
cyWzu+kss2FqcnehcL/Lz3rs/a/bbeR/HBYpAmjx8Dmr5dVVXo9Hn6E8cdnBl0DQFcx7xR6iiBJE
vDQEGibkvTc968VL34K1j62LuQbDRPhk2xvqL0OZold7MGDuIP0G4lR1nt7bGWe53TvAb6BzGhGG
VHhgkra4XHrBweSjLjlJY82GswA2YlRkdjKdECldOGkwzRYpm5xhCd6/QhEU2MD+3E4zjOxxVLTA
+Tpeg9zl7rCNMoSPYUAuS9X27oRfKGaOPS14rvq4WxdN0Tm4GvrazrM+GeZcSgtT+jWdvhqlIAgP
MuS/42oZURh7uWauTjKVmXhic5AOXbu3jsBRm7HGFXTLTprYUbP4T5bFk1SMPyWQpQosMUcavD7V
1r8kCEzOMydwajs+vBdW+h8zN73NgLdFJlsnrBK4U6hKqGUsv+dxL1m5KCxhBhKKyXiDBS0kJyJB
BSIanwzdYSnfBed+V7GLvaSyowhmbnx3cPTOBLETlMMefkaQLvreadFA/qIaMNQ7YdgnEDp1v8nI
7Llcxam/ehfQQIRffWFc+OYMauoJZJM1frbpHzdYV7GVXC8rmlTR3TtelXLYZ2xEm3TdzyTU6MVE
8gxor21zQZolRrhApCyHWBGbjyAolt8Mozfodl/0Ikj6TxXhm9KWxIrZxxf3JusUp74rX1wy7Gyw
bRvAuNNfqHY0ZUIoAyueO9Cyf708Q/0pbXRSrFI8LjOvVhnuyWPvaY/Q9FWGdtrqu82WiE4YMQuk
EouNAbSdRj1tQh3cLx30eaXM4HGC71tzoy+u/8yZi8roIQgXvRdoldkpYViNnp1Q+fjQajZyNWoF
SQC1dDtuIzSFy9JISMGAK61DB5WxnS5oyOckjwuT+kmt/S1fBolYstoq5RMSUFn9yQo+8DuSEYsr
2kCWDIxOemroijDff+4msIL1JoIOajZm2DdEhteHARb/MhMWCeup0gAZkdYFkxcCPKfHd3LQqcjg
EAubNrBzY3CoKzZv3ScbykfO4KFDXaQ88/1zma0SrnyMYEQiS7zBEmyYCXSZy2Xikf4/ryc6MGpK
OQlHLYtzp4yiZfO+DRCjV9zivKttSsgQqmcQWKTG0bI8lZV6/rrk2sn4fi1Ro6kxmgOGfwDSKuAI
lglYXkh65leBvp8sLIwO9RMapVuRRU2Mw0q6U/tVyz1A7QXgE4OWPywLeJ3nRYPx5DXbVYsHAI5y
0blLehpyUZRZtVgbV3avzkSY0fsM3FYZ7aFgUXKfIriMT/KEq1+MKgMnDnlLU6NELPBYSoE+ptgY
8LX+SmtVq3H4eJW+j7LwXccqpM5NFfEFtL/Y4kO+lUw0hxW9loZiLCY17mM3rQFtIyoEVCcLVVJZ
0p+0omeSJijSbf3NrWbqUWUEowCwcSH9HztX0OgyP+yiDUAjFCGOk6vJF5cXmNpswVpjmttLFN1o
RF17Gbxbs8Gtfx4BpTyxDnYntBcenSYuLUKPLtKUhxtGcznMlP6ZpxgqfZvtMAtGCtxwiTZ3wbK3
m6fe0Dxq7Lmf1qzOTWoZUqUqHKqcdU7rsfaDQqFrAiRpaX1NetX/8cyk4PNEufD3wPslMbxGV03/
2NKan3/xQtt1MfStynRiaYDCb3BpWfroq/ax2JrRKuwHygCcVZFUtaDEOC3XkQ4tl/Jy7k+qVstO
MOH8f/G/PbC2ohspsEQ3bV7+mkko/aDPIR2MFw99hP/jGyeKPVIVeYnEhtM0Mv2j4k63hpnzxBFm
QbEDsw3vFyax1o1ZIgu5thP1Fz6j/SIOs6GRHQnm8lOSHtvV8tNeNSUHQOtwk3QxxijtCGbLxZ7L
O00v/f1iCZ2wPzrlRFb6T79Kko3uk4hm1+lAEIW5cQGCA40RLw3OHZB2jGgWbJgjxj024QAYgsTO
HYD07a5L0e5XA3A39Un+d8WT0n4Vj+bHStrvhY9x8/lFZeCL0OEwcnEs3Xc1d7EEPxseoXqcQdxz
/WG4LTmaDcnnht1d5QGhqx2IELw1VOO/7mSinxdORP/CsOwgA8zcX+k1eaBpF+APem+ulLbu0+/G
OiwTxTHAfEiHcu/G/x6zI8j2AjxabJh87CPdvVaAGLblx7+GyjnJkWEvhGNJocIMXyQTRS2yCBXG
oWYcH0skYD2NjTAv6AqXlDIFTOPsiF1WGN9wpzHK5rqX8rfl2mSV3Qi7Pf82Yf7SlpmcSYZ9fB44
cjlOnUY8voC408Aa3Zl7cJL3cANBYLxVEydPfTZGI8i8BwwIeER4FcuGCWzb6E5xDGDy9omaJdST
cIaqomwyguXbASO7fOs/tkwftGRA2fx4a9v+6JqVMXsXqVY2ADGV+0HMkXwU0S9SRXGjsLc9qERw
1WOpgNLZqAXWhjQNprXxyu4PZbKZy0VEIWm92pEmJQEGUdbFYiVHppLfaezZ7ER8AWRGaJqLasKY
UdJx85+U+7Yd+rG3y9TtHiQFIcx/F6pcseWvmDRqC29ZW+/D+98Ww0UaKlhIxengtDbKympnKHEG
fxEjkFI35o6gqdwCWVzXSNmygy0I2zr0O1sHHQpNkaI0OEFqJyDTsAb8zA4wby1zJY0bQqQlkrQn
Z9gpoy92DF6eCOMJdeqp5mT2YifbBsuA9/VZxOBFLT2bSI0kJMsoC14+belMqMXoFr+wi+YU4Edx
r3e0qHXyjpQhynzPmMXVGRrtE29hzS5rqKwqniY22iqYzIhnjECC8nfIyAyoVpFXt9HX1YE555Dd
wUAUE3/efhVBRmd4bngkREhISyaprhUINzVH5xjnzBkJ/B09vdDMGNciQQ9cyyMLXQkfATwDBRQB
SaH4jKjnkJ1l7AAhQDJcn+iL2R0sAwdWd6xw4WOnDd81RyR9REOkzQyMCiv27DWPO3V1NocHjol2
eCCGuCaEkHvt4SmH1OQ1hn2C+EwhkzAEI3Sr06mGZXhYi1EcFDTIhckyew5vxpHfh06rLJyVdmq/
wMlcOF3QVH5dnmN566iqO4ZFKieKxucGM8dRnjEvfqPMzehexuq2F7klfQfRRDNLnC7/PaWHRBHW
PqLFPuW9T2GU0NjLl7e99NXBsF64B3ZJNQID4U943Z9S8KDypp3tTonSizv9tELD3xR6/i8CRkvl
4z/rYzIV/LoRtiek9aavgmEcbmS5DrjLgjBhOmL9EW0gKN8BlQvVk0M6jw/4yvd1YizuUmwrXTad
a8y5clHqkE629Xmrv7ZV3Un0u/0sACuFS9smS1TrjVOagbmn2KnfjYR08OzYGmwcQhd4Xu+M00Ya
v+uQrREnGb0+3C2CjTg/oLJ/sLAUgH1XDDBa7nHtcMjwCyJ9j8n01T+g8yI2bMSa3yOFesGoqGJO
mNcpsnDtBLwsO4/aIMzNqxEeoT5S2fw484vspbsL+Xpr/FIGf2DfG41/bHojlnfYzBOdqYYrs8bO
EY9I2ZeJGZm0J5xMyVAhD5rrdWIEN8KUjKVuxiZuU5mZjVThD4YU89zSADnxkvzLVYAorIENH0UD
cF9YwykcQCgmBPtkmryEl9fc+FRFAPKjPQJTYOHvjGPtOdQraatLYemTB7cFWF5e5eb85pvBfNTu
qr0xz2QoR/rXBS9tMNIk+1b3vUyYWn50bHh4SmwwrNUrM0hILKs3K3PfY0WyQ48kWAFqO/bik7yO
QO8fsnvFJyLzjVyWDMgrG2e7r5Kxgjv4m+iyO9Cd6SyWiVtFVu35B5oKpmwHavkWW8oS+rJuGKDG
l3zOn1Qu52a25jsGN8a4c73pOqvKsxSVKhmAXFY6wq3rhAbif9oMxZQxYFtrqn/irybXVcg335j8
QIH4KnM/BmnCwpsejS85jsRRE7kNxs1BQuiJ0fbqUB+XonDIbXE3yqo+BaytrgT5ZYwAqdKWtWW7
VaBAqFxIX+AhXA0+XVvEzAzTW6kUeBMJjGAFQeLSqnNxcYN4869XaN4p8vXYIoXi/KDew1l2ygrE
5BtlILvsYPIlop8siAuB1LHcq5xZT+5VvlGkXrKd/F0AOtdOACycEAFNNuZzENRVYRBmMYJR3nKQ
TL76reAi/GN984zTLRU3+ZS7EqD6/WuTNRQXaA+oSrkgjtXFDX8PrL0mVk4FNGPKkapUt/TyepvG
7vai+ns1kIniRlfWz3HVnXDULqnxXm8eTcISTbZxDfoTAm41fsWGXOxRd+UJ+TKSSvQXyQ5CwORp
/amWdPre7ZIr3eJQXswksaWFhPnGwnoutCMZjhL5S5j36MD94UQJNgBLncbiU0ec7sxtB/QV5IWD
LtwQpi6mfKjJLRyx8pcliouAY5br5wG3VrR7tiBd06W9GGb6DHUbKC3Bc/HYtHsNSkIFGk3y717R
km/fzHUSvlQ+4TmhBVMG/GoESugVB7AcP94DBROjdrx4jcresREvslgHmIk5xr/BrJgZRBWUAZ1y
D+VogguUHNCftfd2CFD/aFlgf35lcTWN1ZEr6sBZH3c6Rvg/HqKgBcqwLH4mlI3Tf4J0dfNuoPsz
uLKSK+IYoFTqkr2Gps+Py/3PuxSBt7O/sdJ+gXm6ic2APMtRjkhOIuniR7iI0LdByjX2K1R2mS0G
htYfS0X2YwUNiXabO74LITwAN5HaMVbuYseMlsQkaYpieaO8k5YfzRHNl2s/V6FGUkECLnISdUV4
6qNBNwjBXLaYH+HmqlYW4JJMKShOr4MPGw01tTF+TZ31BBTaoC0SrEnW2p6lmC06JSnF0k9cPT3r
8Ax89cnx3E/ERMxp2/iyWlnENFwu9UJPxXZFPMUedvW7rZEQ2piAvqJTMlRpfZPm5Lw6ki+rSQXG
jKrYLk9+tpa3PX2UWtY0eO7AN+gT4y/3bPg/ZzmeY1IdMPbQKGMPfytYuu3QSln+pnNzKsfUZc2Z
6ZDFu97reGnxq3DB7cHverlhJjPGTvqPRC5TkhC/gn6g0HtOTDT6wogKhwFSBPf35lObTYXI772k
z61BrXgG9CATJfEeeLAJq+OkWCkZP5vlMoCQ3KEPcrVcbHk0HPMdkjuSgBVdU1w+Z3rgUJhBvfMi
uotPIREcrli77brCVD1X9KOwD5CjoN3SolK1dOj2XaoJfPkBRg+Oh/ZoEm4js7/KmkSwtM+QTJgS
viJxOhu8jit0OfEBhGTRQPLVZG8xuEEYsdOO8tXPrV6i4JFcO1zFbemrS50eFYL2g39eTEwNvZsd
3yVF01Uswi2mfnyAw9o77z71SUdqc6wg94sjz++ZLN3xZaRs/hJdcXz69ZsLdJuSDUs47/4a3Jbp
O4aYXgNgJMZWwASwFQbbW2Fh6wAoc23BAB2rcUUb0ETiMTsenDjm6wSa7YdPybmgecQWxLRtLaVo
39YEU3D5dilyiVwT7yo1qX4u9Q6xtt+wc8Ad0qK3UHWGDZmZyg1dtK71Ol86o3mYvEx1NfCYMToL
NUfICxYlQdNk6lGPnAdwDxRdzW6onhJRT06KaGLrcg6Nfq4sHrIz+GdthxzsI8G2ntlaX5mafz1t
MbD+5D4Rgdpcp0zxHCv40MrkQzlNDUjDTI6TmnABOTwIcvxtm8N0xlvfilLnmMZXoR8G5DEEOpyK
FELIMCUFibLdlZUiGWBAEgFeYYD59V1jChbh2KOPYojYPgNiadARsEiQifmiLv4CMhbJKRIotPoa
ReBmiyl1wJhkWZ8QjKsKITIo6bBf6iBWGju/FlJHVegS0tsKkjp6seS9lvGhM/5AMW6HwmxM4o6n
sgGlLivJEDxQ11glSzJu1eNHjZbRxHcEn573ze6qGalS84XHQ8yYL/aTn5YXd/QuLqyGcaCuthHV
pOcDGjbIpioYV3BhcUVNmw6qgKaVd/UwtNTApq4ettoutVQdU/FpEllJSvyqd61A1FMt09UEXydG
89GuiKyG2bl8LvUzVq8JebGDg468pYsnm2X0F/IFcJgOkhDApp1qHzV8YzweswaFePnq+0Q/yUHJ
cBNC75Vdc8PhjgBjuGNhJakEiEi4VWB66kmi89FKOsCM6x+wTlSiE2yfncrmNSmHHsKCgrkjPbD4
SMRlgd7n0simzVe0WBYvf9AG+XTkhh1Dja5J68MMr0l8se7Vvr7OhxXD/EdFDIVq0ZX8xUgab35V
LmWTXS6LEMfQt46rlIsq9ZiLNXTlDjug1XMtr1o5v67I7BAoSmMesSKHnHikS1JtljkFF792RemW
uB3T+FvbH+dM6hVp5P/gWftd2VtRO1NMMWMn1cz+wJyvYoYMwj3H/VlHG7H1xLvYQTZNU12hvOtc
Pmz7cdMX73I0NO9r+j8CFlNdP2avyECAATXPlAWeiZX6Q9bBZVTi75OBvKJhc8kLZCza5zaged4j
3NvLVGsAgYfeluRxfoVuyDbJ9hDKAR8NC/pDFKMnRRomJYwcmWRz4X1tICgYZKUqiMmtK/VWK7VW
an6stTAlyy72BUaiG71M7OpaAbZXYxaR1P7rOqyecsoZg3zmsgMwV0GLJAxpHZolM6aSyiat5b3G
XyOD3JOwLLZki7VkMrxq3vGe4kq6wuqLwyT9/v6vXV59IonQSRnFqBuFGEvx8QMrMv+kPM/Bm9uK
suqGrmTkaqUdj36r5pVvSi3yzuIjh+rEZ7LjUXGytkhv8VkguAhfGGRtMpwrjkQL366bjwg3gHi2
CL2uroiWoperCHlV0t1C2Bq4AoradIGa2xzcQmbvPZxLd0+sG5a51qqujW0jFKtwB5Xkv1Ax98f9
roqGnk7Olv+eZSkjABRZau43U0uFxlkW+Vv5LJg399nPa7Hk0C+uMXI3H2sRoXOKa49iiT61ZCRT
pVRGdBkW69gEQOZTzVqniBkRWxX0JHQ4rNiyvu+Tkm6SXdoudgVND5KC1i45LjH2cIlbxsrF+IEP
KXtxPpnRsiKTOz/x4aQziFzpzojvjj7AaC5XMLt5sRqP7Lwo3jOYK5zVhvKyU5L6TXMmwl5MaAnt
PDD3Qr2P7pQo/rSuubVmQu2MUJHodReAmXjwOelW+O+vOUk9lw2HqFDPSj20bO71QiEm+p6QYjAU
l10wz2Sol5u26HwV/paBMshSeSH0ExtMvG+WC6Zql/peVKpIk80yjAMCNf3PyEQZf3JB0PM0yL9A
reUGcoaoMpiMPh4xJYAPKVtXJGmpyJxMw/lqPuBY4ET/d6eyOZF5SlquVwiFwUgkzT7UnVmMuIQX
gJtm2EgepCxJxa9TjI1PXJWEJYP1KUGbRo92XqoOrL4g8yQNOtcTMLIHyD8LkWs/s8zaoZoMOWDU
IoSLq8rbGYUrBgypzsI89CR6XdbqFn0ehMsv1GiTQpb4FTIdFE0+CSniGN9DEy4xA2Z8lk5o/4oW
asSvHXeVvxNo3aAkjFcn65DiF6WJPLeMsV+Z5Q+RB01OpYQ1C0MNHMIekIP24ylKnkRr/8RS/lno
8CXkBLlt2isK5nG7YCMexAvdd00uMiVwkXfBx4hsN5g7o/ODVs6thiAkKFqxJTSu1O3XcjGyMP7o
XTWJU/vL52dpK73aJEBiShOWWsEYAbLbM57TqQgd8LvxUlFkvWtqyLhMejFZUBuapumfsO2M2F+A
ZBsJGhsels3izL7r6ykFhtP/D0mYyYbZbLrn6dWU+E2AxGigbnDm6HKbUI7OFIfkAjwa9bY4ek0f
POAnBiS2KKVbUjK0o+tLHcHPDM+F4k0sZu8orby95h9ij4vVmZwk3BbFBA/i83h6k8vdTNau1srU
SEGleYPtUbNW/N3AqqmgWsgGjFUjF27r+bAwErXcq5RbncsZ3F2bzCtQe4Uw1pdHtz4z1tHukvJt
pGeyP/xWFwIKIhP6fEsFBh8m9vT17LKQMfo7qYz2Ye0sgG6rI0NVoyIaz9StHHyW0g7InY+xVcNI
DkWRrRNqgLhcHXmz0Vmim6R6Puft35XkZ5q9/ty6lDsjZZ05U6/l59dVts2mOLlbNVqp6qmAPP9z
AZIYs4WhJfUigcBWfnhpb42OMTF+fQaDe3WxZYdLnsd+M/fhT0unSnprjDgxdEPjD38Mn7gExgyB
Br5fpEoE9oQ/QjAdbUGDjV7Stsx44xqTJbUBKykCK+BqF3R06IZoJ4MBen5jqnz0hn6UKLOvBBzD
/kMMaVp09O9DysZaqy1DIrmv5i8N47OEiGsFqDxGOMXmdERq6IWji1w94qYuq5/H/fAJBUYED9DB
2VMfD6ReqMyNTz2AeX7meljgagr+mPnnrGJsZ9y+m21l/ETdun3KcCEU6gebPEDnHQCAiupbCNWP
GDPeuCpNDt8QtXRe47u0Hr2MlZ3jwM0qiQHx8udbt8kBAAJL3jQTc+Ur4W10YarFnEzjCGYJu/9M
RCR41v430lp+XFYhoK7CR+iQcYA3/4ygqMRQO38oSZMK64Luo39DiIFVkFjEccsyMtTBkxCUEvN4
I/5PmFVry9wb1/dJhd98bX0aD+kR/tQk0J8GLip++8vhJ4G/WVKDxEbq/ACXBS8Co7BwBn4g17Eb
KpBupn41FIU/Ms3RnbJPlf6tOra5Ay4h6PIMngPxNBghUAbyc6bORG+jM9bnN8O1gtkYGiP/C6na
wQ4BeZub5/1MiJLxT1LdIt8oL6WffFqniMsucPch2ttByeQ418qyWJceXehKVB/8IbpBk3tkdQ7B
hKEbIMLW/XaaduleXmKCgSTVTw0gnUO2I8M5XOHcVbAjfY/pxb8DiJK4A7ECpNoIMqySR88aE9d7
dsUWVsDLuOotFsjXbGoE4Zt+1O8wL6uCOxTbcwLFv54UqCcqu+KSk/bAfLdSILnczP28CyOWuVMY
4TOSIVgE+DNfBBldtkkP6jIeqsNAVTYG2TfNDxXwK2y/aush6NUShd5hqOne2qVluKkhX8FlrE4f
1FyWy3fOugpnzmbxG5Gol8yDIg0vvdzc3KcXuTwkmGXzFg3BmHeRHLTMVjsfn0V9HLH11oDaoVTA
vSJLGHVssDs63rBT1k/x5WGE0Frg1KSpnzExryFqCDJ4dJWLbqgDqzIuQG0O5fg0DRtLHbUQndjT
PMeoYni0hYt4siGbRNpAm4RmZHkEl0dtFPkFZki7UgnmXbdlM5VbFSsv4YWL6YmxDRCw2Ish0fDP
nAx62DFWMV37nqWZJTPSxjKLSbKWY6bRvb75opULX+YbiLopXWgScHLwHmbfHUmOo6t4e53ftu3X
TCcyWeC/19VSLcZIm9p+PzZu+pE80lbLqEcUwlO39klx1IDN6piGi2AtnJJqN1WGgbmP3TIAgR3Y
BEsVfEPYRBv4izmh8ZruzWnbFMz2lwtCTSvmkZdeECyw19vcvcabeGC6C3ae8nRJD0IgCIQrVbS+
bgru2rGiUY7d0ysCMr9riKq91r1p36df0y0Bk+cMP1JYaCQ2wmAlwBnJ0rh1YxgmuIYMT9gLpzGU
7bXRMxPpLc6cZjD36+UPo5IdW6tkZ+wM29io4hNyV5oiMxvKa2ZXCRlFhJz/up77pNdLhf2G5NT2
QYJCOm82B5l7qX0s73UcYB7z2ETu352bG3sgI7scdqSn6jM1pXnk8/+iwaVUlIEuftZHrIlTkWBm
VvqWAWPHRhQYllgfss5cxi72WEPppf2pb2OZRglQYMWjzk4RbTzq400TXCoiI+8kNaCk9IWz0Emf
xScum+rsl/8se4dohtoUNHHWd4sBhqr/Ui/DZrFF10AN365SRhKP0aH7NZB1kiwvOzTkwUl5R/W+
ktkAZ3ArB+Y7XQoWKh/u/XGVR1Fv1+Hom+sfgOLfg4YyohmDifeZRe0FGC2E99+/mLodAs7RmgPl
pv2XNP4NvnQ/fI57PdckwcywqNhPFyFDbCu3buB6+QzEHIka5H9cMKYwbyhJbqCaFKeU8/f16izV
Y9iHYvfAsi6UISuoKJsFjAtkLk/8Av7hJMNSrNrdaC8/GK0LA1aJ3/WwBkc7c8RbbV61QjX3om9m
DbGK4e8JuIioWksHwlsq8bAxFLZJKgW52SiKm0BT2vAuz0hCJMXXTTAwcgOi/kpVu6oy8tO0nMEF
++yYfvHoWiNjeejt+Zurlv+w9gNea9d5AtPtHMIiDPUfL+eT6LrZNq9o5w6W49RYhpkP4VFXGwAI
/pxYfp0PzNsJEAvBPVvQgxP60OrZDHnuhxOSjagoazlIOAd1l21sWv7lKxTKPVLuucM+E3l9oDB6
AyahncqymMKw2RJRxaZQWpeqQE2rykaxBamxD+10pafdaZmd98dWEuhWnQii1L0fFKiYlhwUGSFp
VWN/Ar27tyW23PS37o7WX8n4U2b1URtqmdqpungzPJfLFI2hYx08AlX8WYpRKyu1HRbHAsCT4gTt
9+5GEj1Uk2YBCg+vdmlYJgXM1V/hpY32sd0arc/AYxxFjhSHHmkx56A7JNgarZwJKQsrwtEJg8fW
GTx2hS5fz1T3K9AbwMilK0vt3MoKnigxaLW9/SHl8Yq7IEUOWVf1lKVP7+IDNPCqQ50a92GJTAxu
+1lxEiaP3w06NQzTE7smncZU9ofeCKCTl/0KH+MdkIPCJ85BJnONbSbMsceQ65bwTgRFbjVmlu/G
p+QGpklHwSgZqnjLBsI64PHKhLpzRrPBl79yvfVzzwkRqjLvenQy9UtwTpOVsoaeFWQYUiQTcpjj
Mc/zveA+DbYUiMG87yQM57eXbLYbwdmBoaZchnWCV95sxDMQgBc5P5TJvd5WOUZOOGvRQezErraL
MsYMuwyBQOe04UOeUbDr2ydiEMCiP8P11CmvHff2hA1yYytjNPQGHm/j+J7I+8/weXLedClK02Ws
uKfRao+Ot7AFFWxHuUqiopLAaP2t8jrMOyQQkECv1ypx+NNNBAxs3j4PjwtHGg0+p1jqaGn0TDXb
DlzjsWiDjXP331FUJG/8vEVuS8CTKc1ZWUaBK4x5N4G5ePbogjLY704Ie/fNBoYzAB2n103ymgG9
AK7qWNqP1VTr2hmV1aEC7cETlon/zmcysrfmvowEWeYY0A3MO9UJVlRYIbKz4qIZE5lyYRA0hDsC
O1ebUYQuif1hKvobvzXJAD/AOeOhJaJVX7qbN0chSyDnCT+4Wt6zLojtvq9Q26mem0HKh/izvbMe
MlrvReExaOca+wbTOA7mpCHoOhd0KA7RaP3J+bQe9+k45aKP8auR7SNfQxpSh1AyyzyUGJ6uXQoX
16xaPKDbmGEtN9JADIgRXMTuIq9tyXlN+S1Kg1wpqxvWmyGGnyReiPdFgL+tzGzvoJUQT7zwh5gE
nOaAWBLSpDm5C3hCLW84XALotLDtNVpS0SVWwlFP0KsTNSYlRHdv3lnlQPHb8f+rFGidOPWHJ+E0
bsMaN6ArkTXDpINSOYiwJxaVIIQ97a8SNp3ECc08G6fNQBagTM8iPWPQPD0ORwj2THUE2Hy/B8Av
YC1sTyBPxZty1d+SC9hw7Vy4M4l+IYMxucw1CPYH2fHuZGg9vghYKvBmMfUVvbzmD+QAe4HHN9B5
Hz59NOCe8kxcHXXvGyAJvjCnPkX/+xL5BibgfWh4JEnZFHv6Xsm5te7sPfijb0FDJJ+yXmYXPaY1
WJhjmthZBd1Hoed0k8jIqqUONS3m/sL5v+gR3raXEXd28z9B6i45myrwAzZoFsh7+lR0jo+H7l72
t61f/zi3B8ZyLEH8P7xyE/5aByFKdHC3gGOk6xYLpGoIy2E+Hhiz35tTy6SnznG9frAUzHZcYMg9
qmLSM5P1UCa0L6wtkBOZGLHbhvVFt4/d5EIv0qvM03mJexd9bRIYa8x7pcz/8NF0PXpd3ysLPJhe
t++tDy8b/sJY9elvFwGDK9Lqy+5cIqJzyBGzbhF1mV9tkldC8gdac2LdlUKQcuqXJ7vc0j5z3c81
jOWM9e4MKJyVdCfqVynZ63vwmuYBuoz2Cdw1N8qNCyCqMtSDkG1EuP9tEtrpb30hPQsOqmMHQTBw
7CrVy9Dj7an8g7RQvv+MIM6+mMm+G4GG+HlL5lvsSebsUnoRuIkNipcNpRWMANqry0oOROgGdiE0
ucKEPgQ2D/rEN93PEI95hs/k60pKGiCWSNyn6LnEpTylLRuLTzJMCzLcZmhFZMDw02xJ7B6xnBFS
vgv6hndiDo3MmehZPibTFXSF1LAbTBvb6fabEy5x3uA5gsXJZYm4nO0q3sBlQzMYtaEr+H0ho5g4
b1C6ZW0kbuD+ELq9zVo+HaL0dhfqhJJMc2RZesS2Pc+lupqiGwvcFfNderteLOR5AkvRM6XznxMH
zY3yvtWBzhK34LW/P5pg4+L0DVz/0CimcjBp8L6vsVgVdoEETI1HcnYeQlB3vXBf+9bqPmDlxGxa
23he9FWvpo5rgepJP3xr2fl+JWSLxsB5uBqs+DS+V0kEH1fjGsSJ+EiMEVU2mfJ/DUO6HNs1BAAO
1W6kVz5987mfHLpmMZ6nfzjBuMxU3f0rYP00DTDAPvkh/9Z3ZNcUkwyYgHA2CJvRph2h3cSU/hBu
tR3MZVlXd03ef3AbA1zkYWQhtiJBmjo7cAOjA1WWA/t8Hyuu48XO0L4ZR+rFZRy4Ow3RvqOCLaHn
ixqDfneeL6967juUXcDWOSvv5P/cXgTSprnkk7H1OyoNaBHo2CCPXDX0hhpkAVXFq4/1vxymru8Q
jdbQsGWpfW9ZY/OaD2OoDZIk4rSPBBMpe4+EP2h8AxCEcMcD2T7JY12cNvr2Zs37pZra8PrdH4AD
4i2trJampJVChyzV8Jy2m5lORj3gvRBOxo/8tt+oTHhhwKegMgqqlbRuwDthjc+9lp70BguoHx32
/rKFJa4U1MHvPeHVEZoTD1qNKbt2KKSnFlEEWnuw/JI0gJ2Uw96duMNA0I+QUgNwg56qc0XvcojA
fx4l5ARN9xvNUIDPtyU+TYjEwz0vrKBPu6dxSaH2pu+blElszpCbOjZ+rlCte6rTx1cv+oxxWL9R
jjtHgKbYDaPcLGSx2lZ/MqUWo6CulI7Ln4RFpwwr4pdz8FsuRtu3dz66oEeQXPAFEtjYpjeGUZMv
oGuYjZGTocT29jm7UkBbz/oppln2gH27g0Dx2E4VmTHZFvWphvKNNUNJoPcgTiW7bG1Wf4c31e75
tnp5c1Wm/76CKfniih7Sr2O5cT00aRiH1A06t8hG3XJfykF2w9o5Hlwe66ZcAjTt0hUZ47dbKk5t
T2jdAF8nSUE1vA4T/2NvvnmPY31EnHB//yNZIc/ExTBeGqQC+qjZlHPoDZYFHmKwY0MWnSFCQEWu
g/nd/FVqkfTmnLAYpIK9+G2uTLpJHh4t2HWn/vE8OgX9ixYqZv41a7v7FLYk1KdiuR5NwaJjIgTp
q4cicGMBOPNK0D0PFynSPDisSSTDBrCRg7/6BdGheK2rIu9QD4CXYyOsWBHa22zeZvr7Gzq5sYxx
ot4XTp/cOZxVdiw6cwRj3mx++QcwLzCExHUZHbxhsH7cnVTQemxN9swuOq2qMq4s8nW1nSN1eKpS
DiruU73bzowB7JiUn4qnsYSTQz7/OIykoFKa1ELqoA777Z9uT4IUVlS6OQLUgru9DTfUbQ6ECtU5
NoAaRvhBId4DqajWbD3Co/766H0/5l3Deq1OjUtR75k4u0ig2lOBW+Augp3ZuxHVYGTTjtJX/ZKm
iobe7RBhPWLHs4RaySl0wVWptJWLdkAcw3DjyMJOzsPq8Tyg0kJFwTt6cw4WDuyaZM1JkQWHrUtO
Qx196aBP4tE0nu7aIK+BaoZ4A7ZAxBIdTWXjjor1bAf1BX9+Dmj+zjo8gTaWhiQ4Sr+oj+RAp+ls
J8+sfGcVBI2T4TBhepTQDiJK6GH+NtjQNVvhdsoKbKrtTBtXI5UmpDCPWFwN8pDwBZfuMLbnMqtJ
uJHmBfDUA4gULdQF7ZyH91Yo2GyglBmx6FjsYCMbQ+8icY4tUSGEaKjcSRy+StOmTcL2PvBx6gBv
NOLlZRSw/3dTq00RyzY+CJive277MA6DDcQS31VuUiuQymop2RAi+n0JYBVCkzp/Tj2QD5G/YHGd
nN8S2fgY4PtZzpayjJXPPqZ8Vep7Nacu0qh6OS7pXSd7nQBeDQLS9OCPuLyrDNiE/eyuowV0LHV/
hK3Vv/nAaf4JKHUSh4lLIv2c7bgV2kB8v7bq8A7R2YerjxNVPh3VlSqua4Mx8nwQlJPtsDHMZKY0
mXcdQr/zFwvHjnqkSf9wecmvcLvXpBa8NPhl8MGMd52jVfQ6ESbgqL8xQEEemP/r/abbah1Zart9
PWBcQKAXNVvWZ3KIOM9kIdT1lyOtHku7Rcf9yvrRvhWDj3iQxkZMseslCiwXQlkfFKlde2/e4JBA
dhlqX8wKL3+qvr87Gfm9ww0XAsvEjIsuVaXD3WboZqiPce14gVPwLPnUq3GX4pFNLmjt+vVuSXLZ
hNQN3UIyFP14QHyN5c/ikexgzstV+Bb3xD13Fhne3rdmgh8pV4OlvEwbYMiyv0+6CQSgq/sSsU4p
wMoINZm1qcO5gAySqqEgMdYXXmvVU3Mg3KT+DWeTXSlqKETjGMBo7uXc9CIdstNaWQWI1dIsdh1F
Oe08k7Fodw2FxmTZMt2ZGxYdLmVs7aipIJaqP6/PGpJ5nHN4wryyPHqicSmRPtdaXFCAzT7aSu4g
mt7BpAH6bLkXDw5p8cGmyCJPrAdQ1NkKLXxFEKvKjG1fE8bgc//aFBsdD899wi5vEKWM+Km36Jt7
Pw20u6HV2rEXpQmgE2zaAzMZdTQe7n0Slp3w5+AC9CWI5fNvhl0RE0VxdhFh6QJK3ujsJ9oi3FUx
q9eVJvSY6HKegqZqZvRfTbwsahS8sSGxQ4U8eYIMXEBYBqPzOIhJU8zusS9lkfC5JE2GB3hkO42r
fhvy5EzgGHFmwFL/Yb1OXqU41WjhyAryX+FjH0ftBjSqx8DCu/Y7tfjNvpU6UqNTmSMNsOTTWp/h
MT574UuIOlJ7ivr5wdWvEOBvpfPBBoVqbvHTuRcJm3j2Tm1RTilKSCx4a+U4QrCvQHatlyuwOS65
68/Kk/v8s61/NNNIpwHUDesC4H4wkR9ZKR/qjEM1XNvwulYkIp27cSWLXw0kWr/ASE+6wRWgEBWl
n2JXAN9p3TqTKNQyGEySeHMWlSvVaUQAkwymFlzp7OmVnQYmJRwp0tuLU/RU26tuI56f+hU4nptZ
MIWOFyg1ETbVhOPqLwTVBhuhzsEAF1njOj372MLxFOQ2QjGWS0wrMICyoBD0OBBxogZ1o10u0B6h
vxPNcyEwf5gklh0Fgy3w748BJbQ3fwdTjANPmAAqfYEfJmEnAPAzmjYae865aXj+ceJu2WrjPrlm
olXoJ61BU8Dpr5ewYDZ+94ZNd8Nk2ZRrxPIQ3ZnutaAMJacYF8srXXYUd9HQq4D+ufCWQhIsSH5u
YtRfVbK7gMdM/hDLyeGzMPAuV2stTR+otWlYT8m/40a8B18MBDzGjubEta9H+77P6hClxv7MVorF
3IMT/XzXgAc+hFQI7nLGguhETd6btQC4PxLbQteBclxgoE8mA7FjqwCnNSsfWUqY7Owh4Uc4EpNj
z+5S8UDdgW8W+A2DoPTLivwZpRv/AMcLCVcs2pccIIUnWmVew0KAvh7Npffa2+5dhC+Q8mc2ogDa
Ye/WM58mdlHgSwUtFx3wCfn9jeZaZtRN4JrDuJ5zA14RjORVYlsV3GMxBwLAjt8ZBDQDBxykTLtc
WJLqxcPUudl7hEgbAsxPD65CDh89sqxaqCAM9bKvr23+hVYHkN/XyuTX5PhUU3wL3XsOih+24QOn
eJ8qLhtr865hu1YChE5BipVN5gfZcGeF0qj05DzetSIuwaN9yBc77jjp2Ld+Sw5e00hIeB7e2xcG
vDqIFn7nGhH1iezeTWIpPBdUgDq+z+7AOkBWRU6M09e4osQvvAd+aBYGsODf4HPA6A39CNvYRoau
FxkwMrkeJxjbrvc43rPC5nJLNlcfS8gFo4ZSotWlhvGPFgxH0Jp/0CapcZTRBHkEiwy/NDK7rQvP
r9a1AoqicgahRT4z8PKeagPShMqPEvQgdeF297Qb7Av4QMUBV/j7At6MWgGzUjSUr95B1+1vvE1v
d1BwWEtfBy3QButIdWXRmcY4N6vzN3nQxcOyWwwgPT/LXofSXu6HmFjwexmiES/esaRMc8m5xUsB
6usb9WTcoUZ53brt4cZ/iQUXQUMjfYMKTrnboAfFXcFtR5e/B1UMdQR9woa5y4ora1ku3YGxQ+56
3rrNLIEcUIRVpbsd5QcfqMXpr0hrj9E6ZPYFU6jmfn8ZNoVZkzJ8Q5q4M9vgoGusV/fp1GHC93lD
hGHfNFRy1SvwAiduaWcSKYLJTlUOBvhudQExvUdym9dCRiK+xT0iv6LTk9uXB9xzHiFu02Md+kHc
zEo2BCqfL6M9FN2nsnVrXmb8lU09v+60S5jUu/AK1CJ4lN0zRPLUfXW34Gx71qwrg8vFhZq2W3G9
rgKWBDf5ENK9kF7nmRgmXjnqhYSI4Ny3ERDRl4zhgSlj7Zu5M+v/RSwG7Qi7odbvNkNiKkk8yGbf
m2F5SljJnppazzhFq2tgsk+UFa19RVfJrTWQ8PULqzgu5Ktk9gMw31ZyxVvEdDA7RIkYh92aCtCz
VC6Fre+yjmW4dcc1NOR5qeZYtNXPJrLo4hTDNn+g3qkezj83yW/T95nAdWvOJ3bpz0vc0R9GZDBY
5Ussip36cL41jZP1i9Pqx0QEwChS+XjHcTxerUSeUDB40p31906ATn5xpHFdyKpX7EjEAuhttlIM
iWZo2wipDwHKgz/YZea5g+/B/FR+c0Jjg1q+b+2mX6P8+jyHpB4dJ/xyrAppLjjj9vtmWlxF9SA+
nOmCG+Xfl+4ZbLQ9jCW+HLt6ZRT1UE6iOg27iiLVpMImArlz2iSVrzYWwqLc6O4wEE6/uSj4dyvC
krzKwrsvfYBjOcsAQdvj31Vt0OeyC7qWPvEt2sM26EYgySgzFnA8SLOPgADKkvK6u4eBRI5zOmA1
Hw+F+soKxqowD21DbD2W6QHNvMd3ZVefA/XziwI40ckinNzk5Kx+FrNg1bdNVOXdlvb+JV2wyqMb
ju5ILZVhts20GBxIR0i4yy56J0awYzHRGZFcdPucd7oWHxo9xJisKPW0KHzA1kP3ONOHECGTnceI
xvnNZKAQ41h7NEWNDYlKkZ5Sn0Px12Uk957CD5xD2ZLEfx8ygVPXKj4MqBSzju0iLIhY7w4txhXA
koTdUwypoPnv7IF6fY6zHqgUeFDwwat4hmoC0OY0ISkGourcJ+7G6vgspfbjzwUT8GQkmOJFzN2k
PoKjM9fNtNq/vIBxS9L8tkmq0NwXS9V4ESESEnbLmoi4+HqbTu8i58WMQCqpAj35k+6yBNTwDfxo
bJ9ZZHij/8mwnW8+3yNabNaHFhduFFWofYE7mBrP+zxwzrP0Y3caXjK1syvkguqcl44DWDilE9Ip
8bvQ09qjK8nkvmDZCLugo2uOnE1/Nc6iqrEnJVrAYrwrVpRSt33lLfKAhDIfQnZM/+uwlBk0Fl6t
lR0Mcf7wHB7QwNM4agdzqmRvu+RDHuFEyNH8A9PMj4o/0rDWMqgOoVAt/n2yTkZao/iEuDU+AhL7
Vy0lAdvo7rjwkOlkXb2XKL4IvwZoeIEYapQn7YDxQu+frCO01fQbRkhWon1LBR8enHm0IaOFTbIg
YBESbKpbQMMUoClocuTc2b1bDLrtTdMJxYLW/qokwhFaRXIsJal3SrxQCjmt7hMzBuOBSGxueYZh
3pcrby8r6SBRW9ZzlCoihnCc8gpSROmWrjlHGx+jRF0Ll2OzFqG1iI12lrva5/Vm4r5MmgIRGhqc
DgWizcUUTOSnkcmiW07QJL9DV0dEdOJ7VrFUPQGswMpiqFjMvC6k38riw9Yvy6kWgu3q4B3IBVGg
9PaFQkXz6mpzsIStKFDBTW7cJe9x7icjSLLMeaIdwhXG4Wns1jgI9LM1yR5Dx99eKSYhBvG/Y2Ce
5fYfi67D/96XwkrsOBvKdopIgWaAPwEF15Yv2hy/MKR63Lf9mWcMwctEk8DMs9PqUO83Rk58xj+C
a9+kZJZh9t3RomcYVukfPQcUkGlQShihmQNqzjjwgWFSKcZ+uRNlfSFkIN0IOY7rJQYIeDK7hgMK
RUgI04jiLfvM1BNfl1x6u0HWSjvE2pJlq7svxSKSD175K60F5agwKGKzQ/C2FG2cIZLG8uGzAgMX
QG3mMdRo6R9PD9gEqzIHO7Pez9TgyGDuOn36F3t+dYC5lNAUrhb+kivWPXQ18U0IvvppiuzQqGFA
B9Y9dAeS5QkKiBgUfhTKu2aX92bZ4bOvXXMztUb+HUX6OTsz3YRu8MRuoG4NTRn3gSSgeWY12pnP
lpzQQoADgoiY/jzUuRFYeX1yqN3x3jRtXYILwyrDWbZlZr9ceoh9RgTVn0FH1MVWpPGhol5EYbyL
hK/0jhi87EFo6qQlaUEpmvSKWqxsGVdBVBXI45WzwVVzqlJxwRBXLnH98aFLGRu9bKYZD+8baQBq
FwOf+MGI+YrpQAeSE5wYKCo6+iqmKPkMr6oKOUF+z16YLpVu83QuBxQyvg4TV3VBmQtMlbStAzmT
NhFh1QcAv25w/8TrWpnun36gFlbLsJvIn0n+kwGtquqUCKj5zCsV9qGobf/qd/LFwjWXtuQJ/B4q
n965p3hoqQTWcuyWHGITH/lcAWeEOI3hMR2u3CVHvbdX5H1aJuNoRBj0ip6msqq6mEaBJOdHBgTu
QIkvy+2w4aSogCZe7u9wsjUJ/R3TlYEPzn5v7rrVXiD1MeQV4ec+/aUx1Mom4djGt8o/L0po6vGV
rnXX8T+sEYvQFjFIDy0hd15DzKtNiJDSh+Qajnbo6+ezviigxtSaQ5aG+m6L8BxPXZL3Nv8hqUFr
VkUwUH0sQ9XGEsV7xdEdfwgnQHVPKLsFn9GWyrA9iV0luv6LOZsRJLkJ6akBEv8hFuaHB9EeDlY/
CrJTWEx5/+VHIS27ifxmf1niZvCMNR8tb6d687pkg/Qi3z815+Gv/sZJEq+i7Pj2mgrkfLKG7GdC
0J+I2tx1vjSO1N9puGuod8C3yOVM7gX/FuuKZ9tDegr6FmG+AcHfdgtQNaENCm6pc4hJAbpGh/wI
k0mjpUdR9JsqRv0J0/yfn6m5NHteVPtyhVX+8h8RhrYdH3QlJbNrkdo6+h1lUNpHowZrqA6nnVKu
CTzWEsfHd08hOZb1Ye04X8zOKHWeY2z/bFfxLP1gLDkW1xPripHULskaEsN12QCdkExgyqvofEcQ
rHKVJbSDu/2l8xZ8A7j7kri9bAKtGDfIh6Hntr3EQXMGR+OOJE0iBxeNWxM9Izy7rBN+oZ+1xPEY
JBat6f8asM5fSWDAP6w5Jlr6vBbi9lAaXVI9X0XOKILOfaIKiEtI5bxtNUVjLtj9MPQ7BS9+XRZT
onV1Vw9POCP8tYudyL6egz7vr2x38y/xDAHNLjd/s0CdY8u6zgNm7g1jP3YYVer/gCcNugn0ZLPy
/Jf8S8g0/8SQV/ooXwTWSTonpDIG0cFhkebjUeqhyPqvxhb6ETyhWeQUhoeQBj4msoysyU2kdS3q
KzH6ASQGSu74h3MiArUKIXhhUcnPkOFRcg1GuPfQqN74/45qa+GeDfy+9dCpONsxLlhpLCDroPHP
W+x/om0bXueghd350gMuUGigq69n5GGHI8XD5JHoKJQ547/HSsvYTlximq2liNVQnS8WlDNBT/8X
1FRJhNyeSAI8za2iR/eX5d9ZYN3twb3nR2h1C8WMsmCjOeRIxnWrHf0dd3Koe5vQciAFguISTTnw
OZvGyG7iFXcbNmON3wDEdrIzjU3LCtg4NZWcM824O/a28n4oZXUYmPKKJg45tEd0UiL+cVHqmM0v
DmicmIqOxbS7qPcCPS8AkiH8Jo9vxZC2SDaE7y8rCf3XDuS7x059smXeiZZEKvP4gqPServECMUh
pfv0k8O0eNhxM8NeBqQjA36jMRpg1lguYNZKqSVsY1j5y5s3C0hWhKT6LlQPAQslha2wM7UGrGiI
ftGp4TU1bBtb8Laglxi/ZrPA+ScHuj7/soxAXRBdHuBV8riUgWt8pf+SC3azPfAo6CyvrI/8side
/lzIHSkaAcJAPmzVqQcvWUzA0k1rnkV5dpG9JtHdU9I6OfD1suJS3N/D9vgT4X7opxSjGq9bdOej
gDAp6k4Lxi33KYrW2HmS69CIUl2WNmaf05xHBT3aciVZ+6cIDJ9rOW8/Asi5KWuBf5/McVBbWBh3
0o+szVfjFkuplwVTkzrYVHIC3CnQCfdLnX10Qte2akyL0N75WvhZT+SyAfJCkQ8n1hzftR9wypn+
M1ZugNjk+tyi3TUvHq+vuCSmudn28X26W3hj1bkqOAmCQY87PIPA8Cw2hsKxRAZJSoDCHoIxXNpA
B/IRwTjVfPuOVXWTu6ev6apAIuoUyH1zm5SMOvLajSMQJPc/wlniZLSOCNlYbFp9PkkH8AeNxFM3
H2ePL/nO5CCASWsH8bxZwTYlt/ITV//SxdIpX+BwEHyQWh8dGQBNEMs3kLtP69deQaMn9sgOQK+n
FmXj6LBs8PEPS904JUa7Une8FwxRA3sT7Db89clxJSln5tvCC/2Ws352Pv/YVGZoSZxByjdB7Q25
zFGZPT/w7VSSQ5+sCZAiurrlzLR31Ea2DE6oaOtScfWBqClg0ZpSG17nqTbh7IxmrJFRYTCOAle/
9WKQK4OJbHJAAr4edPvmEDK3B7Rb7LgaiM3ujPurQSTutssGpt2+7kdh93q+X+50tVuTctidkEyW
rc2973Q6ANHBRhnjUfWKTN+Gb7WzRP0orJ6aSAiBs/bCY/f5K0Et/yNaFr8yaZF8CVjBtBT4AYus
EPvm67d5hC20AuoVjX8yqCe2YyxKFFigG5HzygU8FNis2O21u5MppjMBdK3u7Z4C4MeZqwNKeJ40
r0TqW7yWFW+sqpU2I88gdcGjlQrnWT/jFrHOAnacnziXf3qZff3BYas8qvjqYEHkTYEt0uhTTCH4
1C+P3XWGX+JXGFHjrxqMswmEdPmOFInEgBJIWd0GAzoH6Z7VPzg0LmGmzfvHxkXnD6shAbaszplX
57SQ3gMDWQNLmAqPcyeLPMaoXYWKNITziLisEL0bOIb43qOaIEfukYRfm20GoXurOrECHJKklKPb
+wuT9wR7sRZQY7WW1Z9XP/j8rmO5KbsUec29ugPvdbNG8wqEFEIeEjkbbcwiO93lDBTaQyID/JtJ
2LB1Ibw1fjXKzSKwyloClYNOipMWYLI5BcA9evLgm2/nJ6hugj8KLC0NY5dAT5zwn6oM+PMljSxV
6E38y6bZ+YShhmJiwSZzYBqUSdJC/dVOE64lR6gyu7bJuACwc9vtoD6vNKBDTtlZUaRHfrYbklfH
4EkvnqPg/cBl469eV5W8ufKaWHifX2FBR9sCJi90uxRgZSTDG4bgiG3T6su5jqbggzQCBDVWX2+Z
4mBgNBn58LXKFD+SBWNz1YTXe2gZDwJZ32UC2D5k3CzH++4BaH2TsurV+G2qlxhUIhhDKxt5TlFu
gU9xNcXTxGDH3aNY+iDOBqkUwThLshfqc/5Gi1E3IHm5oA6ToWdjVkan5465ULHsN/lRNICmV3Ah
oLxasW2AW1q7LRjehIU63wzjEyChAzebZP245sLDVSm4PjQCDA+4llsb9D1nzm+yNcsqvS5hb/YP
Kb6xonGySYrkrD/zbpgZfnUK1GdiHCVk+/6hURtXP0AYHM+lWJa9psu4jihUdVdq10kbhDChsOXC
AibT+3x8b8w4S5RUkfckrUPbGATUJcC/opwsEx/jQFTKOZ1Ie+wYF/B02Fb3ETtWQFD8zFODcCNe
vtsmByHT+X2Np7dQSwPj/EFYpUqiEepDEczoFBFxxRMk3BMO2+frJci1BwG4Qz73ziGxjvro7XeM
qzcxHBA9wSuOXRH8S5S6gIpF78vndUilakuCjv151+046P0WzT97rWjELeWgxcKyiBp1Oi+8hq0n
bpV/g1sWJrzJXzBaIfvt6YhaobUe7Au5B6QQKzfb6Kx9npS0vphaOYo/EdROii/3TXXpkEtmEcc9
pJfEHF6nsw9B1UnWPlUeFskMLNhKAhYbbTnglmxs7/zvO2c8bGu42rCkQBm6B9fHAZrkrSGUHct8
pTYjQshd2WWQooJt7EjU2oMdJPfQ8l0vJfS0m43fcxE/ltyWPYyyPcoQKIuK4Nezahimj+/AUUrD
8ZSTlPvWN1n+EqHyQpR0gQeqXmKTQO+V+qUlblDa8Ntmqd7kXwgeryK8vGwUpqEnKlFNwv2SmI5z
voLFLcO04RvdcYVPvOvsUfPdUJ8V68VufDAMOjPMX7rIO0SLIeZXHUH4MXeGa9T7cezp0FH11qVa
kuIOUw1T9dcmFv5ckQ83QZvJmVhlTyNnwibrweO9cIYG3EH8BDfdps8HYLwCc5Dd6JY7t68tkF5C
fEaUIWZ+Z2AZG34IkdmOYoj17sjMBTKfJYZzCDaz3kxh5oVGm/dvQelAPnmE3j8njAlSUh+iBFe8
FJTYQsLuFUebC9dqdRtjnjDbCwwX4IcdM2Ru3lTBda5a+QPk1O1KwwlqsHIHJTmYvJjvHwL6+0AO
WyMlG+WYBvDbhjgTtGLnkHpTi7GYd7AE/WiAmvTYwI9rOIvl52aSK+HPJmbEHv9OEXw6pQ8aQZsv
hUnAQYHx5nehSVzBKbMo7cFoRR25KeAxnB2ImIUqWapy6peyoxLz44cdsSVTeYdtiByLGaY1/4BC
JfabABAY3/yioAY8D4WzvuAxQQSQz8Gl/DpVkSNBcxMp6080028GXbs6Gxo/QD7LFVxxef5B7xq7
3nX4nmdz0aStqcNEVY84+lmMmqKFuiXrLPSe9fAnhR4yYQsFnHqOF4MTmVhyd6fRVJPQZCSNR+pV
1PApQeNcgkNbDVUFYoUiHf5y2iEIb9xhqRqtb09EEBsAiRbbadN+FV7TMiYMlDlSIRboyZdiEQms
zMJJNc2+SG28NMfRL6jhh5pBN4QsdKgVzWAQT4XcykDmyIm09VfS4O7FEQomDasnx3cxb6oDGIkq
XYuidkpvvjqO4JcHjjG2PNomJeNXOiTRQl5LKPrhLv6JjOyO9aWibUDz2Ckd+vnyC5wmKqmJA2hY
d1FBWCHK7qv0+TUrBvzTUVNHzAX8XtC0efJVxpAmcXPZb92LCY/sf2wLN78WnicnUjVxItZY0Kmo
NuhAfI+IByFX8x4So1Oe5IpEpbYCjpdDwLRZ02J3PkRU/BNHI9K8LbYcT+vI2601aD+rPWNG/UZu
9KbHA+2u21gOuXFhi2rKEE6tGDXVnDE0065S1tPDibOoz937pZNNjghuWtGBY5EH9XCYLmwi5E0a
9P9pvkqilYgP8nXbm6YThdhk0XRqUvCZ2eg4OGcms08OK9ju7ABsmtjKIo9SNYTBCFuDkyzeiwsK
dyoKfnmpD8mJ/j8/M83TBtykOSCyhcqPW1xUaHl677SZ+kG6O/ajpUVrZmDbdUz9jKaj/lMaN9mz
pzuzZy+mWLOHa2yPc2K1w8w4RnhLg1nvIq18E7I8/zuoQn/E4LhVZ2290LvtEudzaSCTDyuQqgK1
2H3xutIoQC1PbWEbUWipPZklUKHz94I7LlCwssAhD3KEnFpv4s5pK4I0tEK1We9cNgr2b37G2iLh
Uwekk0CjrfXjcn0Hxo5R8r0X+dUVaAgSQP0pcxaOiKVKQJftwnvbEepb3+pKza6/n4dDVXfdHDEn
i/2aKE4Ue1OXIjEiwcmiRmigLuVnaFG8ZWQ9SXsZdpaC7Vu2l0D3hZYchdvP3NTaZvf9+9T8e6sV
SFEyePOYZ995CKIzAsxnR5GYNBivIUzb9uZen9nHEOu2MV5HdaqfsJtSLgoX+/VYFTZvk6GgIN7x
MIYcupVhwfY+Wj35GrpKit3pSJn+doo6S3xEq9tZK/bMKlUuEcs+skoJbah/toOapiF/mer9SfNq
NwQ13jfWz/WgQDmzWhlPlP/1/KR1WUbxaJOiicZbja7MM2s1I4Shdcp3R9t7TCsahmqMnjKXAzgi
kEhfWNU3g6pr8CYyvZv/rQiJ5gORRXiQu+F4llY12CjyhFfJxibZkBMIIzwDckZkb7pVoQYwpHrQ
IMQ6/DVZrGUrp7kpEXcByZ9okKfQFZgMXICdnmvXoOtfBluSOs9tjfRYpK2JxMDj9W53fNpu75ox
3Kap0gK5T+JFh7twdULI3QjYxM+FImAHYvzINMWkFpOQAJje5oqAzMohn83gOKFlcNQNZ0eCPRrb
C6gMTNiECZGgyNudt9m9GhxqFEGQ005YEZHgCULGuVHxl2yQKwS9KI59Ap0St5mDiZnsIKfieLe0
0W8/oAZdyB3Yyk9Bcmf5E4qaagyeVRFzpcJxGbbd65QOwipjQRqzrURERCslGbGrIe0cOd7ZtmZM
HRRix9QvgNPqNgA/x+CNb2+wBEO9azil234X2tARS9jgJvngBAT1yiMcfwlx3Zi13bSwko0U0ZrE
F57Plaaecwwrh9J1OGCJBIS26mRTPR85a6V1P6K2Li0BzGG9DtCPtyq9CA2LSQhWHTs/VYp3hFdv
k0Yg1N/Txr/SVt9QXpG4eCR8X1ICe5YjCdQXepgAMNm6rwwTCFtN70wZm/irtTB/k4ISb0st8k34
odDaptXSocsS+jQoQIfGRuHI/jcbKYgEKzmulZkkYInfrXFHiZ9njugWheu9j6HkFBSLarmepa0i
d5YGEL8MtiRb4RHDbvT9j8ixE3HQ77h5sYt0fdHLMUGK+/y8v8B0+KSxbBFfyIy8EYnEDM6Jl5Pv
N4dNF7NiKONdmVpN/J7nnbxDk9/Ry3Z9hrZF7n4LwRsaRk7Gba4oN+tOFn19Z4h7j3hMgLqJKOre
CoAN1TTqLpi5yrGsmvrRjugT+IASj9LVEbr487ILsUWhX4rFbuhZ0Kdo1zBli+hVDLuUALTvk8+I
5bHF0FUMN4WX9+plPdY4C2+9tqsF1V+N0igBfaNDW8Bqyy4dImVgelkqDSfcj1gtf737OoApsgPS
sksu5W5jbDDxlBwndip4/ERabWCavRXre7fzoPygeyR7c1n6/QpFjeIyyQ2RNmHjwVBJcd8ShYdh
jDiEOKCYtQPv+0JihwnhpBqBF1GK1/RCzSmbNq1uQl1y9tq7U9tEa6dbp1NTZW19D29pXkT7tUl3
hS2Nw5NXKhfgIqT9KtMBh/w67U+a1ExL986k5e/Dxb3gANKRLd595K183PYigFKPIFNSmXCQYids
bTY9UL9BRLZEHLGHdjCSA8EgE1J6tkxlXZ/PaaKKiKqVIUlvbr1nTSaTGcg+6gCA9Li4zgPex/EA
qjWZDia1+3t7W3MXzdv/uuWZFzaphNErGAJd0vxVwx8rY6dTbJ5oOWpyW7NHJGAFwqubLVwaklhq
hXzcal7ccL67gkfQuLGSb8w6vy6ufUXVmL879niIYFjmPh+bXbN5NP7H+tyA4BCOP2AOI7iYbqdu
303HX6WBQhEjWUohd2AzYUn5pj9ZKJTr27VcLDTrdKFvV54nuI3WwVTCKdhvmCe/EUCxMp3Ho4Kw
SzfuCJufIWu3RMH6iBBPqmVjX5m0QJrq9x3DwAXnW6Izr4Eb/7RMc5HXUELjlrH/UDCjy5AMbnNg
/fuZia7f+TRuit2F9ZcIOz+IhLNu+/NDya+lg9awJ34l+PCugA90Zs7S3lmT8qxho5QrghASC1qT
yTBnh0SbNolgpXa316Nz4ffq6bTOtJ1cQF2ERG0HpD7/Mk4okyhNJfIQDcw/fQKnoonYBgKKIEra
1BrgeAetKgIjM9IvXRd0m4BLZdhQ1+vhnSiGoFvH28yU3c8mfIyGCWDAtstJVgC/bDnUcfn5klp3
fDKrJz10vp5zlGna4a10o97PGt1/tuN+wKtmHYcvgo7R2AfPUpGtgUhjt9XDH6m3zHqgVtWXARkz
U/WBoOGXIsprMAXIK5IB7I2/pYSB/AUbB5DTkBTzPXrn3ctVxCR2KKb+Bxiro5izSctxYPN+Cd6p
kFe1U+zNVYH/4MYlo0PLv7VyhXaIpKNAqM2JH5LwB441q2DTBzGQJ2yBYhh7ejAWt3CWF1SkQ5JH
E2RZ4VLU04lPN8ng/I6dF55AHSry0RhtazwFtgnys2ZBRgdasAMNpDjibc3U0CYHngGPgn1SB3FV
PyN7JpWTwtNstz1BEVT4bU/AetZTu0Egum9z6/dM44jbcJi912+0LZqiUrmjjQ5Ab1R6sVrNEzyC
7NNf9jmAeGohEPOoEvpE1cZA4FTGfwuVozMqiygsos+6EYS+ioB256X3XoubZBVnJXS/EU1wOIvw
Jl0IkXIXR2AuTLUQHicfmOs3LAgo9FLrNLyO1w8spXA3AvTF2i+bPfNvnP69khd873ZQuiNTFWqm
5QDggY+gg/X4WD16fhlFMBySgfGv8M4J8+3hYsvL0pbDss/0nxz6vxi/BPO+jN9+tjd3DPqFPGIQ
pZsvI+umNw04f6aY3/UR6wiBW3aD2C8xEauLVuswl88K6ugIzAwG4NrXz3NXMc3qGaX65qNqdZ7T
GCw5n8pzOH8RPfEfjv+VjP9I0STvXgkkehJNhIfBfE65hp3DKUsnsjOBUod4tafrgvoMlbWIpja3
Of9PKdiDZyf/DWKWTNqd6uKhe8vGwIp0ncK4Ej51aX23722GBsxK09k/gnhDwtyYhEeZ0ycqG4K3
jgbuPCeFKsbz1UJrGyZFPgPh5VGKBTQci/u8hHQkACb0WIVzOmcp+dz5tU16WD7qp5vKXByv2ckt
Xx83xEVnbRUpwQPRthIpjkWF0eESM5TZIOKkzCqIjR/E7/o2ihtcuwBDUo5zVVLeaL3LR5jT6LB4
d/TR94hoK7lzckTVlO4nTvalc3fsLSUX8g3FFKzV6fkWhKlRsjY3OyStHD1u1GfmDEGZrmBmW7Vp
hVAaG/OugoPAYd+jKjlZXqECC+Xql349cPrZhqDiGyEpxB0c5u0HHFWbtyu6Nf97V4gfKTk9SezB
c/9MtRaRNEc/reQXqAtbbSOsly1ZwFeD/72xAhKXFTWWEXNlYibdXHS2NrLOiyGXLCL7C9nZv+Ww
q1Qw8S1b2EnteZKCy7u7KZRxITg6339bXXqBD7DQH0lMyXLmh+yhCVb0g5xbSNjDEnJxKYJTZTE+
gjdJoEq9wm+ZCPI6kcWHcUS7d1pUnkhH3eNj7X1DI/Hxu1YDRIlp8OP0OJQHHmFk6j3ZysJ+VbPv
xb7MCIDvbJls+5iG2rOwzlAIQ1XXqStbpDtgSCYu/1BPApHCmO/T62iIzIIim+EzidT5UB+0Xz81
VcdiW28FjNNbkZmPkO1b3JUjWg68fyh2QFQwGwHen5b9WqM6gdC9PGXuR8J9pOalYF8bBLNUJ/Ln
tWobszbGSCgR2dF0CI6E5NVesbNytX26FhoDYEH4apvly3+OnqFWARsszKkRvfrdY0hICmgE/NWS
OHWD6OY3BEWdMFPuZMqENlZAhgrZbKozFN+TvvDGhkdxpwHYagq/k1abShknfpKN3H8gTHWlojtg
LgbCBClucnS9PyzPp7S/eji6vQp7I+PeE2TwSlTnhwipxztwTjtheCp/YUnWjVwttPFOwdfnNw+j
EDxq+ivFKvVZ5gENrCp3PhGqMCN/BQdORgw2cuOzyJqXLFubCHmjTjW0AgX6NFAIBhbsSufrbw7x
vNmvkqquB/WTQXiyuB0+/RLlFdZP2DAZlTD1QfiJ6Gt2/1QEh0UZg33wX0Jr5AdZ9h7qTzHTKxbI
mdA9TIg+3pbud/Q2+A5hKyiLXq1Pg+pF8P+ZMkybrB1mPoPGfP67OVua3uXbULhU2hq3FARvLrr/
yDwQqAi8+YJdRBFM+S4vGlkCd96EUEMQEO7AzaeuJgL3VIlu8y9pTmHFB6sKsMxJcuNuJN9HJciv
IbFvhDzCipx4FpufP3F0L4vKmJSzF+0W+em1zL4oaiT/xO0Gedh4/RlljIUdkDCNi8q4vNpYOwHZ
ZjlK3f5VULzvWBV3q/P5gnBLJU+mhfixI+ss+3nbOWIQ/x7my5nxdE0AhsSRe5vrYjsF1By2IvZR
u9KAG6XeZXFIIwz0ZHaul7FP0VbuCSvRWPewsyjQhZPlLwXjBaEsUVMM3q7wVbVCXPpV0v7rR1Zg
HZRS11rVw8d1VHLgP/puxcUwSU/uHAgJd2QJd2jXKX5fQPeXfw81zDRVFc+ZOG4a8gEsshf8ew4S
ZLql2cz8rKVkuE1jjpKcj+tQd87BWf45qIuwCgiI8+Avy3uEb0UIyMF2bv4C5DVs4StDnHdTrgDn
kLO6T/TviBEwDSOg2JZwqwWMvDdcDCpC+i7YgWkKWoFQ0X2SCgTGTlHX7PgNHr0yhhGjFhNp4kDZ
mdousGnCh8b4WuZd4arLPkHXn1U4czx7fpYWNqjrJvwqL9Cv/cWMnvW8OjwkBw2DnpvbTfd4mCGw
+PsMS4Lrj6aO96x1OtPh2e/ZxahW/fdCVeSc7c5fP1HUld9QHWTde4JJxtUxUQnCZBIXzXVmq8Oi
kcYtCXE8wO7x2A6MJJPMuiE5OZBGh+JoM7FMoUesqRcgN8nH4p58nnTMrRoxtBsw9qxcQzZyMIve
g/31XKrqgqBT32HFfYzDbDxHkmpN9emKbVRmeFqWU4TfCAWcl9msxGsf9sQZQG4PqxYrpiGc014o
wm51jLSwXOLgx7LLNzDQrOkupqiqjmY0UIZbD6jbma8yNfDnqpcEcaVEnw+I1wbyqU2kEvT3Kghq
oZCvcKRuqyqHBjNMTWDkDrr8mCqQ6pTb58HsvWs4YHwtMvOITM2h7+AO7p14FRfZvB951RodJsxS
5z7wuCmrOiYkVGs+xEAUJ0JunPMisR8HLTqCgZYJ/PKxlX618Z3Y/ycEqzkZkALI67CR7jXSSpbu
sdgfsvFvPkZOh7dZKcV1I3a5n6weP5Y7hdbtvI3SSVjUHxJwSO1c3SkdxJ/mWAaKsnG5QnQo8DtO
1BPwluHK+ltLmlUwMiKhpdO265Ys6oYQgttm3v98xbt+ayNpd3cx1k7GHpFQt/TQrkDwWYzNAb2/
nDvuWUNpTYQtyAcWu+i4vZcU5U7o/EvGi7Awt1Eld01GDzUKVe26QklgITZDwEL+K0SbDoRNA+uZ
oQnSCCWdcz2HSigeOY0wdj8eQGI5HmzNRMuWDn0rEH1f2vgSEezAYMmYsvptZf5x0Ox57dHnvaBP
9CkWbqw+b+x+f0PC1+mo3bqeEGRzkVK9LUjjcy6rEHUUIIys9bgUFMZOfotMPx1jE01uQPLppW51
ht3YspoAJ9fKafvCbWZIlwdswTw3jk89O/IgZqUbQz6XgF8xqYxCV3LIGdN73Ci7cDHr/rfUMpaw
CVlcdiPMRakXlhaYDl3IArIIiRsR3ESA0jbsI3ghcG4klTVl9BIigrNn3V0pu5rZl51l+yrTuAzk
Qrp6Frq1VhKaqt87UE53kkXnoDYqEBTQNg/ys0KMSgYZvq3shLK/htbva1vgbHeHyekpIEQPmDUE
5wW7s/bTKKZ4eKsI6l6+XX12MMn/dCkloQyZtiGnNavUDKwOVg9wIXtutygOMeXEtjULSBRXUqMo
lCIW75vGbWOmi6e5qsojX3XtqVyI46nw4j1Grlb9E3jKwLYWRrRUPCKAYhJ4hyfBZFKzfy5rqIWh
BSYPaLF7W9N/xj1Q5+4zHTKc3J4JDG+OZ4nopHrIq2r2G/3byCxfbV08Z7e8anUinYkpS++fuse4
ecZwichwTOdL334NdBTMY+6jh6L5mi5U4/Bpv1MveNDVGr9cOLSTDqmjs+8b/FYcl2OEwO/p8Lc6
KwuBIFsHuEE8wKs+UIxdVgAl4mIZ9PqmH7Use94GnT8MRxdthuMCpgF5bRnbRdAIF0fSuMd6Q+FJ
KiZlicWVm1PyInz+EnrrNNo/GLMwCB5is+JT0uuLNlcjBpkTGEwiSKKR/NOKwfGa/WIl/MLKDrSd
8Sru5b15wiMqduy5BdqfaXWiWKYHQcAzy8WdN0cm4lywzgCZo6Kz3m8ZJsTdL87P6x+hGJjb3D9j
8F1E/oC1Hx9EhKBXfgVSGHs9bnBT73oQMg7Iky8mNBlYbrcBW4aU2pwZxIYY59Eew4hNrk+wm3Da
PoafTbW530LPOopgUIEcrptI7LNMXqTcB/fqh+P+JHrpoGQpG8fsmi0beAf4YdRyumJKIW5HoVd6
BpQRuow1/Pl/46JWBhZZshigwBXEaibc9otUXcL8LDRg4Gzjuccr4x0/nCW3VaD+5ewybDdOTYp7
Be1CY8oZUYn6kCGjihxs3sEdCqisyBa2oo/o/Wgn8seKEhsyBGNb86jxbf9B5j/z4LCjrf/4OSfq
VV1ZWHFAgQ4w8gqc9U61YJjujFWQCsNyZjQ3NN/bYeyDoMBTEIsZZloL0CIlyUrg6YOqKDCafL5t
QxzBpYaKV0a9ULVYqdijzfODn9xanLsFoFrGWlJX22CR29RFz/NLnlFDnHyyBUx9B+JSlkb3kBHR
F6g1NA5FBVYG45zB3pkqd48jFQ60TjbsDqJj9QHyY1ps2Qu1a1TGnZIXElS4YJNA9/fTrHJTWfMQ
ZlkuoqCXmlWDjt+Pd+OVW90KaPwaZinSp1xDTfb2ErL4IH7ANahu8vncOYj4xJ1sHYw7b8ZCoQoG
Ix3PC8XIojX/jXTJVdFB+gD6xvM63gAmoUIl8fxJ4nkU6jGsGMB0Z8Jig1g6K+ChghCMGf2fDfoy
bSdd37FyIAM7EXS2MKDTsq3Z9HOoxg+aPnkCgfdqUX/qZf4iviyrvnkMg5hfNUIRC+aNe445cguE
IrJ9qcpn4+DRJag4IXYDg4S2w8bvJT+yWZ8Y91YsCMCOOc6iWWkj+fGUUpGBgBm9VV/ydelFRPqh
s1morknzLZl7C+vDImr4IGqLTR1WOwHCi0oatoH04KqcRm4jUzkaXNAsgsSvdgoZ5Y4ZjLwQxlj2
J2TRv/REPrj9qGPDkgS056BpILP7vi49qH/8tBLuCirTvbpxR8EJ2zG5IwSMzWLXLTEdQwfxh7AY
xnd5Jr/f1hF1r5WYwQ17S0Lw1UKZePzGZuA8olLvZIu/cn3QG0KJ6O8rWmUea7ySjacaU3sybDho
agmRaHWoFo+5boGfM0SN1fsT6X/agzEVRn+rk2vAbV3si2/xFtbD4ckpLvV1Qr+0Cn80sbS3i+p2
K4F3PBpczwRASWZp8Kr5qlJtFm4Rrj9rT7AWClmr1tWPTpNo70LQrg7wR1pCfGr5/8jCAk7r7Z/T
kURf9jC5iiZvc+ecXzcYK2l4yrkzgG2QGJTTd4+xYK2YXo4n87/Z2xhkBsphShoX05AntoO7CQxf
kEjinamlNKVGEXpMlUbWVlu1v0clV+NAXGZmtQdflwJdZijwHJRwhiH37MEXVmBl1kV4CbhrTnN3
Ysww2Qof+WZdmS3PiL/UvhILOJenNp8LvrL2bM0FXsrOG78EuHzf0NuvaJ4c6229HjT7LF9yO578
DD6ss63A84xPzVEbPiSYH2bK1nT0U0VXLRGzPKOgnS1kAppj/LTZsIkoaizEU2gmySfKQ+u0Mt36
RP+zNzTdTsxT0C5FZec1bwAfVDkJkmk3SBO7WKa5DKU+vahZDnnQ7yN3xGqfRSBHFsmM4yDkPFX0
HGzH5B28SbYd5Ztkzd9Esl/35W9TicUxTEVwqEW1gNrUszreBRy2jgmO4Okq3URm53oUkllOazEQ
oji0zYaEfZWB0t9C6Y+E7/3NMllv/Os76632FzDyhLy/sleVxUFuJ9V4kIZj1XuBXPhQij20aqLF
cRDq5pTv5m+yu530C5uqQnjvxqFlzEsC2q1WdZUN+AzH6hiU5EwKkP9bx+UHI4bDH+tZtjVBm+yZ
f6/6wm+hFVz73B27bNNZhm8WCILSFqmPoA7o3rKnaWUab3rreiaXP4mEDQX8VrfJI9a1eJHWKn5T
HGhzxlTPw6Ya7cMsbvF5UIeBblMXFkxnON26L6J8poCWtHIVLJuRhwwRyc0mseTYBa4oNCVCK+Cc
BWapgE1AgNkcuUo5476NlZaIcTospRCZ01GgrubNGjJJ0Bbaz411SfFyV/5gFNWb2dWabKSX+tdn
+JisWXncd/nVxwpfWvSSveI7mHdCweIUidUeOaszyTLl6WnLqNSmSZnAI04/PbOy7uHr4+S7rTGQ
xQo2xIFNjm6nbfCoC9w0YXaZLTUStVVSH2vrbkm74M7xnPFjZSo2/HyObPzwJ8fxoWUxzrkEPc9s
J1E2L0fpEnnLZLfvlwHmkFwlZ6psAB0ZVee/lx6CjGus2NCTNlB2zVvX9zuQaaiPvzQfue9xMxVo
2qbUPcTCAQEdTdhf/ONRsEWDuSh49FBymzwofI0DzMsBwdMlvGMTCPqb9IwIlFtkLcQ6+MWQ73KN
K1woY6phCWjauMJJes6UTpsaIEB3yiylxGsSBg4pMR6v/OJv3dBC5YPJ4BDKS8vwLzcMXOTV1rfG
D3IM894XB53xPd+VK4iQ2z/fEhN89d/eVes8NsM4E43Le1FW1X6uI9zNbxCcLToBggpyQ2iVXdJX
aCkMdivhsvnowshCXMzVnFS2WobOaHzy4RbGTo9GY4YODUUXMMiC4XERgAkocMpLEF+1wvrmRbGV
AbrusUuPaVAO9AIGa02kdpa+oSYczfInnnv9qvg7QiPvV0GeDHXZWWd7xEDmEVcve6OK+iHX02Bx
nI+ZD1LCoC+sQwWb0kbfXwZ3nhEdXo4exPR3HGveLkqo8og91HD7MdFM3iUCj7a6RgzOmn+pcUf8
GeLq3ooNI9tnVd+PEmcpurRyLiNLz540EgL0m9lCkv+iWyGZQxyJhhYsdzEQMacMhy2cE3/25KWb
Tt9DvJj2Wd2jJhLH2tDxwi4qugwczpMIuGYEBz1E1F1ajJq1/9NnkZGlXDd4umLQQpppQ4vgvz66
7IvvQRXpmgidnuOvrIK5/VcdKfyfxm2GVJQMFjKtELtU52csaH6axD5tOlKc3M3G+mP2g8qzRxGt
nqpS7YYUmaWyjBBEVgdg2M8Pr0/fg3g9WdVilg+QYV4JJVjp9cq5ybzlLjdqks0zzWXa7wZCGsLe
ifG1fCADCs0uUfNIMC+A0/EwPEjHtpQ95g7DT76glc0KaMdCs6FAW/JqWlGKywwMrBYhcBPVSSqs
B5NGPxQ+sjart47HpN2+KudNtTUcrzB0s655+ctZslqQNRiQqA4OLgVPPZxX3dYZD723r63cTEJm
IIjlYE7kYDfl1LsVyQ4fcZ+Yi5c4Amai0iG+DRFHRqrtGTJrae0AuqLSLEAbAELYCnPGjUInE7lT
74VzXWtvVU2GO2fGKubCtgukqsBKorf1HWk16AVSpmkO5ioElkGRGz299OP/W+QAAOZmSsANJf6N
RF2AyWrs/ro4VGyjiRelnFCONEIxjIA0nLzigu9+D5nQZIf06kIro36YHMXLdoY4gHA9NaMCrRf/
q8MevtvBoEOuoWQBcJxbooY4OwgdiSP9T3t8BFj1ZBJdPkPMsazqrB3sPH+yFTgeuzAgPkqKjEN3
IMJMVV30SRGfXx/gDseldCuAWN9G73ujnAQHZT17zmsYBss626Q3y5xuH+2MBSrbpWD4+G6B1+MW
TcrwKRnlzqlQyUPJ5qjAUZ1U9De7o2oDS+DtGzR8rjxGSX0bb5bTTF3BZ29sv+cYiMhJ2hKAyhKB
hryFRAh/fbrDtKMYhgA9B8Bc2IoxCYvVLV0RwjZIK2HXmieJGF6cIFGMoEFO2N1hZ+LX2v4MLeME
9J9OK31iUB19OtjptorsTNPQ1D3em4DZvT3XibvRX/WSH8/RDvg+APbLGZnlPWIWeXzRv5Ec+Y00
LlABC3EqZP86rDXACvIWkA2YV9yEW+lZW1Bzm42TWDwI4YhJAJaesdvf0rN0m2UGhGbdY8l3ygfe
cDPBmrrNQRjnXxY6nqvUzKskhrzZrPeeDEuReCvcFQ2SqGjwzt69Aebrfpxq2zWxAzfAcYcMnZvI
zrG7818frPHJXE1Iepop0mRqU2C8S4ytxzdn4IJm5mymFcVIaV/nszUzXLq8L1TPG6iVY3owfN+b
n63dVrnYLjai+EXIMRWYtCCYFNWAaUVdVRsq5kM1xOJ6OA0ZGou46b5pnVASznAtq2MZeR78TIA1
hng3OXzPjSd6wfHuhs0OuxReJJ27scMvhWHBedGqbIXWQiWXkfWiAg1YPEZMFAD/IWdNfbm5lb2A
BjdRX2uggMs6QxxERDg02lxME0Wbc0JmcOowYDHWZj+dEwm9Ql9mBG1lOdHC5Ix20p7SmEjGAFHy
xExk3upPA1Ytm1td6bL/u1ZuPxZZ3eFOuAXtaq7GVLSoQxEcBiLyVutxu+T3zzd/TRcn3jB1DGAY
tfcHSzduq7sN8++kQ8K3WXoDH+akzIhbhCDIrXa4buWiUzKYMxUaedwfrt/4+5wYsMm73Iq8ltxj
DEr6WfLbdispIZxWRnlqn4t/54cECIR5dGxAWW+mFfE0JQeqYfXwTnG+7XWdhLu5RGyJaik85Esg
G3CTAtmLUyltnhyb00FcuWEwGgXYZQ/QzkfwaQgdX0b3qU0Zkhg1fCW9JkMuPPkUrJYf+8e1Iqh+
Krs3YNQkifwPNoakU2Kn+E5iZPr8Ke2R91zaEzx1OMJftUnbHkRm/x9qWLuetkfCh75nSkaFkSBW
/4dmNbu3MZL6n1v7AfYnPFBDy2+dbmryrWnXCshjJMOCbnDCdDt1LKLlpazr62dJd0nZJEM4PnBs
ZuLtVo7hNoHXgMXuJGrpFSmzA5FgfOo1j4+Tf8rfCAu8xVFYzUeuUNJW4bIwN1TQOvGluPuUSLYS
pOKILlymIidpF8M05hMGC8ks8S8oN3bGN/ZM3ECqapwpThPWIjYxl4GS+olKY0AbT7SaACeEs5N+
wd8soM57Ra2DnVQrZIN5zQ+PUmqHSrI856mYr6/ECmiu380qiR0qs54sdSyGphJ5s2255OGjXajN
+3AxReBB8R5vh5mZzH6IOqJPcBs2S8Y9d7HhZKkmnU0jMQT1a8KwT8YH+Opgs0tel5ulunl4CuSB
72/UNSrOTxtbiKIMJVWYGk6ycn9kOpes5yaQoYzFvHXKxedGaS0MmOyuttOSfE6gq6DfogJuMf+Y
kzdg1VGzhRxSRiFNtCQYMiH5Wyhpz3DBMWInrZ41tuOqRvbQYRiowEdU4HnkZcKS2lhflufOC+lR
8yh7pzOWqkIN9Oc1Te/qOvhZq1tY96I815boSLKwpxDCxRxczYGlBLGtASA4JdAJFu5h14tUJO3y
f2FMy2iawS0C4SD4L2KG53ttYWA+ftgg0miT7D2qI+20VNw/eByer8J5QjO5WCO9LI392GKkUYkV
m48B0KplpPBTlEoIur87TIavr/p7Di6nvnVn4WnwPU7NjaYMT7dTKkqQoTvsHec0TPPqCpmoE57Q
kSd5FvZxYiiNz+20fkmC0jatw8maPmSmL0eFEEs4MZ0wfYLqMV5pJu3hCYRO4VCpbTb49u+2dyXF
FpxdIe8G0qBvRS/uKNkNUIKOOA6mnxq9+O5l7xEzpi37mvTltbO2BP2nR0BlVdyihVAvhErzn0uu
Kp27tPaTj/bHvnvn4LuReJNEgXBZbRqAQstCk1hpPL2kowR0ZQnGSR3O9lnLhmcmzpLaGQ3SmRkC
hiGQAWoO/QmXhgd0MclZF4y1zt1L9oYKmaCgqfpQdH6HeSbn8r6O0+8tLV18p/Ug13bUYb/sk5Rw
qCzo3JFQZgNif2wUWLO3UGGcDRo5VEBn3TZ3VDWipUPIDt7H+1p1iQyCLMp9VHKKqt1CyaVqJph1
mDxJS4EDLVH03y1pc5vLQ6i8hlGHvPC1Ex5YSKW5CDI7a773QQS7wCZiSSzgXsyyK+k0r1m/HvF+
rh2YiUkXx34+o9CuMPs46fh8WkFngmmhlWodnx7e0wAjmsj3AgwGkVvmZ+GRjzOxfmVmN/+MIKhl
ow9TRv3alPFiHKYlERSQomBibY4wVzg03CB89aSqE5wGi5v7wnXbO7v66bk8o5jRUtwTJd0KYqrs
uig2HAlCfzXTHls/iX5H0L6RHa1BPfzAml/998lT9hMdwLW6ZzAvZ26Rlwn/17ozpHEoHIT1xu/D
JeQ9kN9EMZg3sMUwCPJpCPHiVkT3dyeOIYrM392JJRzWPSzTbhb2kt53UF0/SP2bPLHMAzfCamFO
UlzVUCa5Hhi9Y0qN6EmI4n4IQPZtzRVBBANus8OBO9pPgs7kqQRP3SWRhkFUxFx7t40DMFT0eRs3
jGMlhwqU4oMVybhZcHO9FZ8oEA2dLa+P05V9OOOOw0f9v/N+oNrlMiBFBQ/+5LzsdJHvyjdXPxvv
LlZU0xKbDv60xtGlK/yJZE38JP4KneTu/FyePu6TtEfHM1EP0AoaZt9SgReByQeC91J/w9tobrDr
DXj1v6ovD8z/1Wzp6KZOonOiNxTH/cdXAIrbyWWVVSBlikpQRx1GmbQ0mZktRzVfhuuJOvJp+nIu
ADMRak4QJ6MZ5Z8qO4mvZwYFdEVTjmWKoI8b0Rtx1JVDeFze9hH0qT+coovkv31Ph6eibSYss2oW
q7CMGSjtedTxOGxQfwtGWYsqCeDXQ0x4p+/3+7tDPIGr7LkDCvG8ia9qlvVqXk7Nhj91fHPcr0nN
Cy6+tbM+6BzykumzMsj6cDrHUtLqVNCNnuzyrTkztUbpgDr6yGYA9Xcx2KyGA2RJ3ccyWRtu15DD
CVcCDGh81Vgj7m+1n6+lIY3417rVP4TVk31659zdgpa6UFKwGZcQfCKSk6JNUj7E2fLiQD5qvwgP
KJgYzvE7oNTqlBqh2La3f9aFECYFomkA05zF2X0uUYKMoLNVFjje9hBRIJgRoNUNXhvBoQBLjJ2V
IPWECGYCl6PT8Gqg+J/zNcjfNB46dJkh+OWvKBGMiphNhl/jLO8LxZLPJCKihKJv0jQEzqWQy3BX
5bmlipfcR13fKgeGlHiMfclWN+RCEfiERXxuLEqDJUxKV8n7SI56gWuPyrzWnoF3QaowQ2woev6B
DOzJePq45NVC/1JV174D82Zevw7rUwEZGZm5XTwWBriZq3vavNbalAKtMOuimZEZVrfl4P6eUJT/
JFivHzufQTx9LLqQXkTiCexLLif9yQp0/tAqcKggFdoLkzbSnj/2uNBG0e3r9+4gvC5EKJDx38Fj
KDuS9SKeEBugNE1DZYlfsT+rSNO0f3aFS5p9JnIilfv1SRbunVUqpoEq6Brn7aTIx4uc/b8CdRQw
ISdy8br/Z7/0z72NWm+X5jCeXQXEnADWgRK2n1zQN9TgCIvzv+tDw+lqj39EkSWvpD0cxG21XH1W
Rt0X6TjAjAjYvx9DV2UVrrqCk2gK1t2lkDLuSSkeubSXNiJzMKTdJQkHU6v8dt8nZIzP1bsc4yCQ
qccRbG9J7MU63fEW/qiw/5wo9jh0diFFUAymS76NxiLCki3+6nHmAdQ3HJUi2y/9U2byN9ssvIKL
ajalaQyVUU0iSalhqobn2Ykg5INunVNn6+pR6mDSb14NLwvwymP2Ty+gFcNNpVjP/xOshdURCKYa
piLF/tTMpg68tUw1woqdM2FrLNUHgcFfMHEY/30SHpzWFMYTwRLCRqF+Xto/at/ezfWBa59gPe07
f6AJO5mMPTy6Hoe8dJkiZfT+uvfU2+OWa91YcaCKlXxVAdg/hwzU67xmMQ37xwr7B+hTdR4Fwpow
T0ZGNgpVn9DlDSDgZoJAUH/Eq/iGp7umSVmaNWU7ksigJg1NSdyDEL4KXFAm/fv5xxZkTFtaEHot
s3myzCoQW2cidHDwqYBzUAudLKH6xbyg9O2/Ag7ZpGMJ4/AbNNYX7Pm01baN5jlxV2xWT0ggSemP
jL7ybJk/P1bhNaFhq8AFlb9uI+FcgUjPBhudlygT4cyxdC6AsSI3phocrCyWM6Pdtq9MBomN7+2R
121jyAzk8zrNQPcA3T5UmFX7QIH1BTP1Fpp1aaBjm6xSzVDuyF+LothKyHkug/ONO9if7kP9Avhb
YmgoQjvEaleTO+DVTT7KdLvEAdc9XRw/sqQi0rD1K6sPJql4raiFEuKPkmmHSgZDi0U8SEZy9hK5
3Xup+uZckeSvo1W1ryCZBNnbFC3yymr4LV4OA2uNjoMUowCApTJFWiho32ddL7YROfbIaKf/QqlC
jdaH45LZR2UOKL6+HfXJ+mwac2DorEnTXUCVNQOs74asw/0JX+imBl+jFm59FdoNLH4A7ExZPl2y
Bpw3EE0JbkbLI+UanYcCAoHPPqrWg3kbu019lqMK3X+6P5hhG6Xg9eyu9xSGzZpOh6zq0oV+WvVz
u0x26fHmIb4lpuK1XcdhzN+8n25EO7g3pKd1PYTpMwoXjBRXGgVeYdWDsGPsoSlcRk6P6nRFwva4
0QzMz1WtVook/fHPyJ4fyqfek1Pwax1hU0J4dS6ujalKQCgtmuzxEFGyKl221JBaR47+fFiOQ2HL
pnSBdqNFXb5Ed/GT4lVzezJAqlrAXrtzlinzqqcmRSW/asF8FAv7k86eZnjKJXvGmsHxaxbGhH1Z
JiB2Vc/C7TM0s8Zm6Z7xM0ENkYO1XeT2M0qhc3BdzgjInufmaZ/QokrXZw3ULPJ6NevqiYYmReKD
IGqWhM7LHXdKISuXiZzG9XLQPP0oJ+LQbCO0hRilfrA9YXfC4W5lwfbIheSRL5bi0YHznggthDWQ
s950cdZiTKyo9pHStwdpYgKl3pEh+wSD+FY4ZSlfRIRn3tve8IcO222llru7E9YazSOJ2n7fi5i4
zizO8jGco9ARS24UX0ysNXVWyWa6NiK/PrToZ8FmxTSh+TKOl1EHU7wNW/Y3gXldTh/HLZZR1bxX
d9jhTdcGoCH1zBB6vZjwVRyp2p4mB61xD+3m6PPrLallEnKH6YEp+Ht0POyITzNW3zJ2akbb/NYI
KybjU18NQ4TCCsUVSIPNwt0ShQ6DoSu7Fa3BTIHUt5IezbJvfxxfDpQR4f7OtZV1Q4aClFh6Pu/I
mCXU+VsQH3SiYF1WWBT0baVCUDDKhhmkn/2f+g2GN0SOs7BJg63t66KdpHKZcwptcZdId+8/xUxF
/9J1t60HvoHmWD46dKHD+eQwqZcRoAyoPV3Az8CYbaji6nwEVN3nnz3iidQ0pUK79TyY/FcTyFJz
oXm/rr2mDZV5ljIQd9sa/0UoHwMRvlsNd2ekyGmtBqpKpFEWYeOoeOzD55qqncFZvnweEz9IJAsb
rQHg6vpYUW3zYnZfuEG4zKV1xXlGlcDKy7jlDw4ZEnuzzdENuUt91M3fuKbSCH0Yoy8eTUkmIhlL
Rn0eS8iCb0RbPfFjP1t5i34fjuoCZvZi2877Rg5r1EOonItUSC40Qacf4ggposGu8OR5szqgDXsL
BfdQtWMU2PJTfI5RpClb8mu8cQDq4F9FRXD6pSxD8qA/l+i4bQzsA+h52Q3P5rIJQSKTCc8O5Cld
qqwkzYYHncseTeeKPyzREtNyP4DHtjMpQZ7r53sMn+INwLWbLNdB34Oq8qdBfhJwjAVexDecQLnH
IiPTbJPgNejFoljGxtXEJbQnblptOtC4KV173JgnFMinz8eZpe1XUE85PJP7jwccNCG3RmUBE6ea
77FtwDKWjs/yNVgdJ/RlpExjkrK9EOKPhMm2ZXyi/sptiVhWl5PtfG7CiLQ3v4MXAogIC6nZ1D0Y
w9EC4uY3usVvTryhoySPnziOU8j90UP5XlriPYr7ycf7a57DuuA/Gxi84vX0btZUzLb7x5Axtrma
NxLy6qpsOMobDY4nEZMIekudG/zdRIzWttzYwEVusAq/N1o2UTUkGrH+bwC/XC6EjSIYtRdceiw3
bDuKnNeloetvPFWGsttfANca8zAp8V2yTnlTzqSTl7KBD3y3JnX+ULasyD2/XSB/Zyje/Jo6Vfel
higrbxgMW9ykkpfS7CUIStHb3rl60xUdjDxK1AcBBSAdJjKjg2V/vqQfh1GBwsjS4ee+FLTdMP8V
jkFK1uapeTJmt9AsR86In2z8zNNBh/Trz1sZp5v31OXTO8it9iTrZ2eaUVKd7B5UcSBPOH8itm6z
ch5LkUkYVTQmQvPnsBKT17G9Ee2g5zg5vGGUeQr7Z/qCrtIAauy16IdFaaOZUIVQDJZsa+Sose+r
ebeuqc6VFYq0aMvvnFFvWfh9QbONvrsz5Rv9+ANtyJfHT6BPueMfLmHuIOJNGLVZzN3uUXhbILlG
k5m2rwkJdypoc8NJ3LFdNgLVSeZv6d/2xmo78XHK1kvXIAnDTmGW4YKGSOTd7n7r+R8u3z9OPgNV
Vs1yYu9md+bdxT4TdskeO5hHXxibWoyhiqrGyKABRVV24YzIbTnwfY9NMvDiw28xY10Fd7TN+CI7
wh1sRbl1bypdrjZdn8CeLViMf12Y4e0cRiRhQaabTEMZywtDmjbjJuVjNx5Lftmtdn38rSG5qczZ
upHpMSGkh3YnDjD6HkJjPnKPMfVciRcJMUFdYSl3EkBVl9PEKa5RoCd4ezw4tZl/DQyi/9f4x2Z3
Dw1pLd8i3pOGi4SEI94Cf7jrMqccRgilSwD1ngIS1uLLqghiIu4jEnQh4X7dlbwXwTnuUGPF9VrN
5tJikySXRaDw0KAJxbvuK4tGwsrdNgckTAyXJfSvb1Mco5o3P82owp8iOTiQhqVfnKyBq7EHzLRs
wZFU3HDV0nPhJBnzOSGbXBXYVDmep6VJnF78vwue/Kvoq2QXND1ijTRjnYEqONrKFfeNSZzH3qeB
nUV6auBVSnaWK1MD7pPR8tZg0hzPPn+MuqJS8nrMS69KCNr2EwUIyZhqfTr18rwWLxqfjIn49maW
5qYjnkGUjekzMU6/jbJ7iUsRVPUYt+HNOnrTu2iMG6Fb1oBF/I03UsE7vNFrZUJanDnuJh9VIlbh
RSCENu9o7jpRrxP2VYbILpq3uBQQv2aSmCYutR7K0D2BrtnSLnnZsBzbxBiSC0d25cI1tgMTFkyc
YR6AanyJbNuQiRfTyE3l98r4Xrj7qF/MVl8A0EWM6m/JZnDO00+zKGqXTgTj2oOOUmeXxyvBQ54Q
ymToPIAtyhbtmHWZFnyFOiWbt26WWbpNJZrNWgk7u5l8Ytogd9JQQpaFULCybB66q4oUdTwJhBgu
QrydVCnKy8RdVDy86qNiHEqW3WLbNm/NBF9b59C02qiKa2YzyCN2bYjGnBfoG84j7jQICA2HFhj7
moj9emqzUQCKSCvg77KHWHp5Penpqr+nnkKbTeg7snO0wjKQ/5xUxA07uLgow1J6Tz1TL4OtZbqV
ptdbZpcoBvRQzghmc002As+yBxPxxyWxp7Um+llakmpIf2ZMVReggmiW7ndfhLe4+/3o7zL24rAm
byTlA7EPi3ry/W9Ov5s+XjNNaDen5oG2MtngeiJSC3MmaG6SxnjjBIdIG9IiBOpdeQc+GurEkvus
MbPzJ0BtDP1/AKWtY1cern4gsvnjsmHOe6gh9JmTNSVMX48zIAvyHhh8Elv+nRa2rx7xOfYr6WF8
E6MB6KqicVDZymHmcmNw3TrKDPcjNBYgD3d1iayWa9Llo5eeaxLdT/CfpOMAfkYhhp0ReJNUkcWK
IMsDSkYceKxjz33ziDKhVJ8bpMP3YE8ONJ58yc9Mjmekrc5OI5ojpgIRr+5KLQ5Tvh2V6IxWgav8
ZzSEuWfuVw4tXFnaIiJzYpBim0TseQ+MMQGocKnTwhm1sMZsFIqDcp5jINv4Jreb4od2ftI3dgnD
691SrcQBawS0BjZVJb5hPgkDDoZTBQPH0uBTa27ii4P95KW1OGW2RuQe4C1udGXl4fo720Hdsw/0
rSkL6m+hA8CA+4fb2Lg99sufN14UQBdFMfpmETpjUQmaJpYdtrweuBr38pe18hctTa/MPwxbo6tR
wOu1k0K2fOSHF6+d9sK298yEe+ng22RF3QFrLD9MQYnHcJr/a+dQ9zicZugdNjHB8O7OnijDLke/
A3LG6iXlF9nvCqDamYcgz4Bw+QcipJ+TSNrabXtKHEbbuj9Ew5c6gVmQTWJHnTZI6Q3f3r+LtPLf
/JtBGH5nUDSU9UCAtnyt7PD9XmWp7NlHF4eEMBeI0V3HNF4q8Foo34CNnA3NppkKczV1pdHs6tn+
slj7Hthvzf+gaOjZKAJaUZMXlqxywD9v763PvUpqIgSH530Wtf+96Zr7A79k4sqsu59r9aVYL88r
3jMt6Wd1Y42MumP/Wqfv7NZGAddHQ+l/PKHZZ+1b6v39SsPVQiiHdoAxB1I4X0XxwIuclOTTP8Tf
frE9Ai0DvEDv8SCDfzaovb+awgqRa5DleqcivzYzORj/98ASR6DWmUQbPSI8ndot1cgsy8W3BZfl
2PLG0xS4Fo8C+Cq+lNIcWW28ltLljKteJpU97hUuMMX2owbHc7O6oXuz68SlerH6SzZLCPeTlP0H
1+3Yf3BCL7FqYkVbBLuzG6V37v0bh+4KzDxOOQUAahhcsatBpeZeHhq/HX/S+gvSBdNrBHGRax+5
9N8CKddzxRHdDzXi+qfkcM1qDYyt1B25/w0xIdm3yMeX4GxY3VDyAsilrAmG4A/JWzcSdaY6BWii
pb1vtPkcroU5asW+DaGOBTzEE2uhJ3luTZPclm9NUrgOJJA5eItAQXUyd5xYBBpecsMU7zJxMKYC
qw2BdVh2jbVVTCEHkTmbEKvTiCyqPx1KZGbpgO56hJmcZjrf6diyiXeQnfHCTx0RwMPnpsh2hQJX
1SrobqpA52NRrH47/n/unBaAoD8UVPzbVYNNpIegED7zzOCM3vfriPLFt19ZYqnxLsXEYu2Y9whW
52WJikgdXwwJsg8WR36aJCILzOYcIFW9nA7KCGbqRRKrMM/DE6fm9KKVIzy3afvhP9F8yDGT22LU
qmCWqAX+tOit300kc7gmQZvx+LGkGhbNb94FzfohMIMif6MKJCvqRpActm1h4f4xK0QKFI71UBsW
UMZATYlMMBh4DZkz3u1zYQJIsGOQmhbJYDA1fshO19TOh0SRfYUcux/Vr2pL5HXJKWVg9pFuctIW
4/MBRV4n/3N3Sg4ZB3MWa6/DIOgJVFMD0ttPxlBGxT8wzJJNh63Sj1/NNswDJqK/7qoo68K/fhPA
jB5OPlT3mF4wm4RedxRrl/xqDmxa529QopNyx4PAPir5ZpPS8YDRQ+2m5rAp0kCsmQrCjwxXLvNV
AuNfbpgox2Ewp3K63bH/8rjLS4JPMuB4HrD6KcoB3LxAZn2eUbcG/WdSSX2NgUbM/O7pkXOVtGzv
g6O9vxT6+eZinqMTi082raT01HBpVtrVvArJUsj5tAjjbm8Peu4j4ZhHPFiMf3BVbgXh/JP4NczI
Zo/UHitwpMvtl/XoLzAlLYmYQvVUu69An3klEAFt/qXrJhsGrwDRuSoEPRE+3U6ZKbvvO3f86/Oz
UmMR1cqoE+vupsXz4zXy5so1G7HFpCFBXUU6OSZMbgfQ+9rrfdPH+4XHBDe2MRZMx6ACdGuQ1YR4
C1xByPUtQ4ygD9asi/OLSQglYI6f5ltifqfV8qbFbxZ2r/brvMyVcEr1kWD8xuAtw0Ultyg8ecdp
xiNncJOq8dvrtlVMKFJyQ/Yfk4Zu3ypPKmG5rZaOKpTs+hp8p33a6L9rTxyuayAxi5tZ0qAB0I1T
wX+gAWfKghthfUjyc55fa5xodBGCTuVaZ8ojkr0Hz59eApeDZG90LAqpwRRkZQYFaYAkpipTS6y/
c7OgJokwstfOUGtoZL/NMdQ2J/dsLxg4tMkquctCpV2v9kUjkr1+LEu7t64zF5h1m1crf7R+NuLo
3WzBBUOhuqRCR6DWnUDG0I36aFud0O6f5YI01nYhrcszpVLb7Jby4FqPJHMNJBuoWTevkh48k/lJ
Xn5kyD2E9pWdMNp3L5pkg+rO8SpIlFxrfburHyWc4Cxe0m6dvg/nHCU+j2oJexClpS8JEGqgBa4w
amNJ14Oa1sTo9jnyY4tTIFirB0TmnhbIMxp9VIjaJgaBTyJz6DM3Ga8Th9VSaJfkRjDh1FHszvxW
OffaIXjZwEl/BJbKulZ/ihVAtc0/fmRk9O2ew1fIZpEbzq4hV0KW//a5sewJI/yD1EOIQHZGbyFM
6d3zkJvDkpblFgsQc5KjEVkJZJDy6n0RF0GqaNZ8MLOXcuqaAcbknojtUpqF51exFxNi6ZrIJyWF
hetdGVH86Y7jj9UfCEhv+Go4Qtsfg7BpdxF7kCGTPreFs0XEJoHa9sJBtnIKxrahR+MdwmhFsUY1
LspztG3Eh7V837KC3Uexu4CeDNzY2vNMHdJ8mulBh1eDpQjxV3SWy5VHSWGiKE4P1lquXmI/lOE8
40V4nSf7haGYRW17cdLBjMeP2WYuyQBKbd/f0LPHVjlt53fDnMTrrfuDrZYx8DoWTKdUEbSRgPs8
XuzFZidQxgI54E0sNCzsp9VUvV4K4Wa+mVdyAfmPo1NlX7kjbUsdz1bgqyBG9Hi/vzW3ffwmepJL
a2AkESUP2NPeECtOa84Zm3+h6VcDdrURp3QTR/hLqj+vD7SwxZVRhJIj8IV9dwY50SRSwWe2WWgg
TxJjR9q4o06r2Yb0UboPvIk3hRA6S+EAWKPsKG06Q3I7FHncDYQR4zTAsupMoNM9PsPg/JqiQBna
71v1njWMDYx8VHLROSpOvQauw4A08CYVUbS9aqubAk39xYzq3kgCRnAXmo35Bk5XYgUJ82MwmbHh
6imaosMZDmVkX02DOs0qQTncIr0qnFAL0gDLZeqeAQiaCgKdipSlkSfj2wmAShpeBPWo+JEXS3Tk
s1wX7ll2tlNSFbv3NwXujEy9WjWKA+Hwzo+p7ex9DdZIcAfsE7qW0fOMef2JLEy/qFqX54C0EIxS
GgjsVkiSoTTR/SlzKxxfcfjV2hVM0LDk+BP25euyle85SeyvfPEfEUBc9S8kCEK8XfEOADVM/spX
IdvCk932On/V9PCcu3tDsGuJaq2r3FW1neHwlLaRAFvYx7JcyRmnm+lJnLpU0Qw9dop5roixNsHx
Qbhd5MKR1FmfRNCl3DJSuD4onco5sEe3ksXo8HoHAwGOAL4V4YEeQwaYpcIFTHQj47tJ/Z1XIxrB
ZH/njFy/NkYIvLCNC8HhFSmsfbEa840QujI2xLvzZQajc9g9QK8Qd1lkXRhZEOJ045FvEF6uLpor
Ql7qX3hLEfTlADBmdUKnQGR0UsYKfEpCe/zwB+nv5Hy3EflGO15VLAzHIqBn2ZAGBjnTMCFaT0NO
fdEHAVtQ0iYB+vICdpeKFiGZ+lqrmT574ZN6NlLmCn4Me3g44xO7MKmnM9ShFDVEw+I3yVjbbbz/
ufp0ojJkTWxdNn5gxrQ9PPxj9uD3O5Pdr8E3TlxR0huvvVJXSmJ2KQ+hewPesyf8xhYvyfJweQV0
PjqXvwmvpbwfBj0rfVAxfke5RaGWfP+ugQK5yan91ne8VA+6KPPsEMIo3RounoxRI9S94WA6Snub
uizS5eal/xiqbqDgvDSCiLWkqJidOesbKj0DWdwtDg0cwU1dlTluxgMpRak6gmBrdJoERvkJlLAV
vyrRlDTvDzV3WGsQJzy2Q1XJjta0KxT1KKnZH57LgphsUnM2s+MU61XWspN2TwBGB1C9LJNM1bJx
+tmBC3+TfDjp2D/PiwF1nC2FxMNVRzt99VqOsKuNKe9FpZ2CGoHebGU8GaR9IQqvda5AUk+TMbmI
neiqTr9UNgPa9cfdgKpAEXMFzHqkGaMUxAFDZcYmGjWvUxjMu8BM+/quPShmVrJ+AG/AAGO/tYKv
yWR4yADDMa++9c9GTj1APx0dyJUsf5w4WrYdUEldSgr4XH9F6AzopMH4o4xRU7BtdqY8ey0WDuxA
YWs5LRWBWADr4I6ydMbx33K6x0jXx8Izl/JE44iNS6d/vniPI74eYYKTbWbYf0TD0dN6EGIOBS9c
YNwYQUn+uYnFPcH0QZkxKe/D9vILmpjwMrNk/hG/adqyzaBcE+KJIsx196TE06eccYyyz0NG5NLi
KA2D9wwKGfCrZPp8edPPlPnUsWBU4XMxfb/xNAMKv3E8cFXKw0tJiXrSDVYdXi0PQWrJ3+CFyAnz
2kGSS43u7C3ZSae0VCX1qQrVCpsYfrfYcYaakoZa1LVw8WpCZMKzXB79UAMQBQ/iirfsZfRNd+Bn
rRyjk6ooBjtRBVWvt43pPCKkKP+l/twmZL+bSYgyUGFeOmut7MhEIpOBeeOyyTmjemVTnmXs+E6J
orE45dur/tiWJwNjpwX8OnKe2gcaXYF2UI8uoRvcWMyMLnOSw7mYax2xr+f2e0g7wCdm4UHQd5wk
AYXeEeI9kvLLY0k6A7AT311Z1FVQv/ZqcvVDW4xHDuA8MEu+BWGeMqGWu3XKeDMsZGaeM6fuuie4
zkdMDsU4Zecq/Bq7I7GMbSwBq6ya7NMnn6NS9Z56YWc3KKvLbFWjAlaLVn3kwrKJJFMDCAVNQXz5
CyOveTOvuyOjFBJbp3ACgM5EqV7FqwrdYKW0Jtt5quSvZGXgcwJKRHjVUpGmYC3dOrjyaZvRHUGh
aewjalPobZZTVcPul3jB8NRHDPZx/120+WDqo8ssr2tKxnNAgIM/NgQ9PVToeUlqSTjuFEqp5Dxp
+tdZjfCr5Ql1OzCw1qsW6x5D+zU1E41vKvjfalByHj34mUwZd3LNkCisSE6xZbarVVRbvW2uwwDm
svJ/T33oNGUo7x5RoWNBmP17dmA1hyH3AzBHeErR1sWGnbz2D9ggJIumVOYMgDUqQV23gq4b2PcQ
WXY6f331QwS3vi+JCu0R1RMJf+rcTRuk0LZIgwTGS2vrVUskTEY8llt/YuU5e3ZRomwBs14xRrdZ
7f2b2jF4CHcYMb/eVypYyRgtCvfsaTDGPHs6bofHDohN/EQumxQcJWvyV9Q0BwA8CMrNd1LNH2hf
uNbxO2p7FvwbgienTJQmJybDpjNduUGq+QhDtMIpEhjt3flo66JkU6tHV7OOIAXuSyAuUQCkkmWd
z7QiPw2lWN7KfjUjdxUyh5silH691FUn5meLPBUy6QC6pbk3SU0lvBj3CC1WXbvUuPHLiL/q+Gku
jDvoZOhnakarOOhCrXAieBc5CyV7VLZ3BIcun/cEhwk9bpasBJKh0jf3LTfBoEE50Cm9UckH4ibF
UewRcgqpPIs2iZj+YuVmyoQ2OmtiYbAdteMQfNphSVHuYxCdqrZAulHOjKe3ValNC0Qq7u7dds7E
jXpUmXyAi64fwWit/6pGaLeE1Ib2xvwllIDj7WWnPTFrfpLX1i4x1rbZ60iQilXLZnHR9b1J+uDT
4QyaOlfhMykAj1pic8VoAR4b6zJ8a7sCmTa5/JuNqznyaNs7ONApXrimM+hh2iuMVRYH6NxY03i4
39IkV90TsrcAd+9KtbPqr6n1kGo5WiIQVmEZ/Wc1gIH+vpsFGm9U0GQaaY56kOOxXR8fAlCDHu3Z
3+Li3sNupx1S02oAnEN4USejkykTR7yjcp+K4J+6MmZRxcvvJNFF6YivFhNI/BVO1/c3uLcVaS3x
el+02xyr8v+ZrAiXzqsQpVCc/yYgwNf4CquFkNhj5BM2smSg1iCpV1FUt63LIN4kttFmLL22ZfjJ
kzWDRHbL8fnK5MBiMLhvs+BwqiG90a5BLLuv185YF9LBTdNBThDcyiZpd2w+E1loFrz/ykzrvlw8
xiw4bGhW1igs55r7iCUD67PhFkEfoHPEz8DCgoyoA8bLXts/7LiiQijR8MLgtr5nTha7+BOeSY5L
x5WLJYO5XJywf3qAIOiSVoRHwff4QA5ck6OJ3QQDWLCReslIqhEXnIjnWAGqttXXmKvHgH6kJ53M
xDg2Ctr3F8RMLnF6G8e1IOm1nned7gUfEsfca7e+Q0M4DQ1TnnXjfDdpVOZQ8sRqyOmN5X3yJyWB
tHX7e9xcbnQBZ7QtYP+GmQB9k1eE0WTr9idbA/6SDFEbOvs/NydGAWnIYaNl3hgDsEXqWsIoAGKQ
bgFCiSTXg8azBPdmAk0YtM/GP5r9HwwrdC0rEcFPmHaRJjg8bmyQvDfjy4qiY9CGMCKRcIaThWXN
I+1sE+1LFKhjc0dQjnz22BqAncbIKOxK7DaLpRwsBandkdFCVSA8cSocbFYevg7tYvE3q/QIQpPH
wD21ASiodPyLkKd6cSd7nDVTWeSuCAG9Kslcxi4oBzus3/pzdkFVwJX4mOJhMHthvhh2BGK499Rf
qOjVNCs28f4uUg1w11+HtbEdANYZldOkzrK9xN3ozQpBqXnE6giPJelYVD+D+kZKCVKsM1ui8+De
UnbMy9T1JYAcmvjz2Gxw880srxsrL+bMzfwNDMLpLb5/V0y0PHBR4UlXt+WLoyatCe0AtbtNjc3l
4QV6Rt4+EITeJH40d7xqnUQWtKOUx5se7i2QeNFaFGdcWt01NFL1hxSSCiS75t1n6ua2dE+9G1En
AzFj6ogaT+dNTFmJON8XtarowpaJ7TwmesyWXt8iSIKQ4AzNOflwKYOT/R7pTEU4iU617M6GilRa
OcIIVln6WDcx+lJCiLa/0/F7sPz827eCt+fPaHTq7tjtWenttz1+p68DLTey2unuxYjt9OWO4Zqp
uJawp8lWqJ8L0gESIM/SQht3c2srrs/53nST+pSRC0vHmEW90KSyHYZ4yeZzaNbNKMTb5ThwB/i1
uTuXXMS7b7SQWxyqyrTgKmycBPnzU1O8yT8IZTmwGpgYRA/4oVVfCfri3hHG3yW8lb5yOrmHNstn
tOa3tmoZXiVg22DDvT9haFr6cwofwkYElNFu0ok70KdKEB8Hp3GLKdnUxPPnKa84xceFj2g8Q4pk
ekwFC6ak/U8ksr0yoWqNsF6ZRPXKC2AvnoIhhypp9nWvy9qsxgje6MZ4RseVaCxMtIk8qlXl5x4y
tYJAjimAVTkHlimcagwNSWscJPYcJEWnOARNgHrL6mmOHYYb7p62B4p5MPGJBpgzqDh6tgFbPG95
uDRwOXeW9z4SZk65MPwuBdzOG90kupV2B9R2FK6qYWuRoVeg/ofNp0w2QopL6ojMHt0YNWjdU142
wt4QxbhXUPO5wjNavGDJqo7awlXew+yyHGxZKnE+DB3DY2LnJ5M3PeVD1uIgkuKdpwkwNXXfnmK3
Bg5nMO3u17xRTDSnc/TFK1u3UefkIswoV9mEOVRj/SRtgi5+YGx1819zHVMJ/kxJzet+TMtl3/ic
NHI4zoQdjvgbBs8wHUiy9NPJFb9ZOcPepcXuxRsXrUxXxtZ7sH2FInJfgu+6kHyhpYXK9TTWWhEc
uhKLjgQ8z6s3NPsZDjNUU+dhAIGKkzUR7pQ7Ynh9eNsXUiiFcygBRZl+O+zNf+U/2Y6nXk8jGDTT
MDgcK7+6u4SCy+8sBXeFZO5ZFix522sJ+Nwxko8VLJssWlHOKKKApanGQvq84pImgymGvQdvp75V
yScpRLXpzyIHlXIYKWEyjOJMng3Vkl4J9h2rYuzLpd9ZUtexIjbQxMdmfclBL5GiW+7AF0AqTazu
c9wDpdpkxyrEtUi3ixsv2ga++XCgVt5Glh02rfHn4Ra5xYx7xt5T0L/DylfyALmefSOlSqfdfRKp
m8BBvo8iV8KR56NfjaSeySoi81dc8hy/hKILU5LphogrX6v1jQp7sjfsIwUF4wAlQ4yBVvj25aub
RoJ7xi+TreHli6EXNfEoFELdYY+m33kNahZybRvF4QqafoBbhxxXvq4z5WikW0KmP39diquBdW1o
KVCgL5aSa4Fq/dCCOQHakQHeCtZHH1dosNZub/CSOdIw38fGm5kHZfax8BqI5PEYGBE8Figs1i1m
meyCxn25fc1kGVclUnQmZeXh/bTewSRncjqAhBxdxW0PytxNFWNYEiyPmUH9JqeHEnRfELmBhkZj
IduHrvyBNTGy2QHE+dwpDM41ZYF148/lOuiovYPuwSBvgk4nsylhyCYEAMXhef6EU8GRrN+q27uS
JM2x1JqiIar6D0CweibYNIVuhFpsHAwftiRJPvGgXH6BmIjdC/9qTtk7O3LHuEjtXcwKCVSTNtKo
ObaxiRjrp+v+e11naWPNqEI09J/fpk3h2I/YEfFJVPQqBouDJ55h0DdAuEGJ5WVBxUJbYU5xvM4P
IzR/Yq+EwDPJDg3mHs4JoMdfGohQ0Z2wzwnt48EQFnY/BDEYBmW4NTCmKX8Im56TyNHrzoYt6/AO
tcn1igZoYb5a0Y8oddDfTxoFxrdKsFhuVeTO/GyJiiCdH2G9UTvSwymeow1F329rOnlNEHnOWVPX
A+o9+LxSCfH64c/JpeWSqWJKwbZxT9kXDtmwkz08/5N04w27vOcQF4kjwXKzJiaGEGzDULmScf79
5sM9xKa2ZE2P4hLu3BM6IkcmX5yp+TgXZfdRs6k9k4Pv0CmlHAWVbF9Xf2J/7CpbRoacd5ySmixf
uzhVhfOThd535iPSAWaN2dPgJVae5xf/0Wh0xxw5wI13UECzFZYTAebxiwS2yRsIyPu6Vg0ntSga
6x7jmU84511JAZhKaDvOrslPdGGZeDQGYq9qSpm36WgkfM1klxWqbL4jowrVIxdLj69EjS2DYLu7
PT8EEyU3qcDmP3ZV44IEzRIoyr3zXaDqeaR2E0uPaT2oJmwKKjnRJO2iCDM+JuVn3oq1cD0dngAk
1jcQVG/JQDGXnBj6zqto5ZFFIQkxxNRcsZXSuhmGLurZnctFAanewvZj0JvAo/0OI15w9atxg3Go
P9YVWrDUBDpkGqbcmYnGrq5HoqkfgmhjNXzpBiCCcIB0b/eyGk3zPxmPK9qkFYFVIsgK7voBZmzZ
+M41x18NwVFIwcMX2M8Xf02K4y1cFP1F2QsIIWiPGRF1DjMZjtiW+W690BVXcsSYMWrnyxdSCIw7
GxfKvVK4CCrdeLxCWDfBeblwMP5W9pRvbHrqnDSTDt9cz8NBdoz0F39NLEfqaMseh0Bt4IRKz66B
dRDlAr1PhoD0PJ8i98vLPCef+vCd857hvUOS5JuEuRq+6q7Rg/qc6cuxW4zfxH9mmxHFC9Qv3fY/
QL/q3BZ8DAj3Rc8oyKCf3CNr7lItbDCRIC0aeYvNYCpbs4YW3pTeooGKR2rFFXa+zo5TJb5PvKNd
xsauJO3QaxR+zKhQ4k4UsVYBiMwJQFh+K2Sxq8wH0531Gi6eNDWS9ynTxjSyaOiaoQbCBXn27VG8
E7PjYcXcAZ+m95AD7ke8YUgEyTujH4MvxNWBy8pw8QCwXxFCo50gKvzuzIVP2HPe4s4Oau6kTqVY
r07blXCPrV7YrZQ0MZ3pGWRpQaSiRwgRS1yX/gLB1QO/g9g40g8OFNGb8IB3+KGg/ZpRcJ6f4IXK
nC4GslHKV+SJD5nAmy5i8GFLNAlaW1zQW4wG+F2KiuO+gMUHXQCD8S7t3jjmoAf/yJApJTq/RrUc
gBhniocDoUy9hzZjcc/VAdVQBUx8gmcGCbGr/Pe01Tuf1IXp6wblHhTuSeMHZjQyYjwaaq43Dn09
R6ZDA2jZKqpvHb/qmQqAE1UFks0BNZPPvBzeqw0QeBy293OFOBGSXuL+CcotF5DlJuR0SaIX+fGt
wTaOkKtWsoSmzD6Nrlb914d4+fp1xbHLInlA23xNGvFAMz5W5GzIOxvJvbCPb6pf/LlEL05WPpY2
9UFTg6yyPdKhsK+mfsaGTDLxekkVpd9JdkkKM4YcvMV+NsmOdQ/B1PVfn+4uq1Tf/R4BA17Lm0Te
7JcZkYx06ZA8tch9K41eEFtMsMd0ntFyS0drTZqeTd+qODjWYpu9JmxpIhuiXNGVZ3DZqkw4Abnk
c8b39IWc0XAlAUh6w82IbSnsox1sF+cYoskR5Vvjmx3LbjNkB3lYlLbzrUuerZou/ePae4Y1Q3aM
LZ9eAfJO3T3GEsB8iN5ez/Ajjowjd7mZGXDs8Jb1Ys0FTKG3wMEW8xkVYm7/+OprWC9oDfOSZ3xp
eEY5/3QZqGWpzfrpy/UaIAMtfcvalMq7MdYW68S55OAKfbpkZGur5JuK3SgwgQKKozYgTqmsG7Si
8iTNS1FhMFo97WFmULw+1mB3EYtFoc5VU5Bg1ItoaktzbEwtWSa4Nkre/sA9w8C05yTF5tF9fcWW
n/iGEGKkUcvSbd4Npr8YakXWx2vUBtwzkgLS2Fxou6clS7hn4pILN3UVaiJa+4u8BApeN6oDRtM+
+wHTa/dMm+195p1SG0SoXVSIHrRGfBbaZAkHwsHp+T/hmHHP9F35+1pltLP897WGV3EiB+tYbSqj
pibp/akQSAHqNHYn0DVBtEpSSZKTDfRIevegAQHlNEWOOdVpA5XtSOXJIHX00l3C0LmzTr8zQOUD
ockjjX8KNj7edGjRHQw6fMQ/V9xxPHanfA4Aiv812r1hAg+ZePZehgb2wDfROqRoW0zXMyHnEvrF
U392oJlJYFi0LtdyAdcFlzovBWk16JP4biaqRkBuCQUe7bMGp8em+Ero8Nqq+V82vD4hC/xwwqZi
3Me1oIz5va7Rk3pvZ0lgdrkfYKXC55gcHfPss3CmlChOXkHX4+yZf69314eq1IbfmmHu7Mcq/CJ8
Kg9QtwN87milPJeLP69G3Wch6pcTr+NVy/tYLYT/aHmcM7ca0E3PoRyKHKXQEOWrdiGEHhL3EL3p
DwRvZ7FJawtO2Voq7drzJddgI95xgT4EeOvpfKYzw5RTlYcAjx0rZSVIvNAewIwrSL5OrdvWapWg
0mNIReeZeQwpHDkTXLvtX9YiEOAYv38LH18kZ7Ww1NAQjD29DoSWPaJksuyB8gswRQxQhsto7E3R
/7nHorxVXSBWYFJ5C89uBGRoYUmJJuhCthk2uKDF4RsqBZWb3E4w2TlYegbZUGYAFFAGbPdqHoB7
NtqcwufGVLUxlzN5wiYdoXPkJeIkg9AFDg4Fob27N+fwmA3gW8eWcd+pi36e3YCYIel1NgDQ0iOl
oeilSTN60QFzV/tiKjq+SIsLHb/u5WYlzLCBm0u10G0tmR2W4/SQi5I9cJSvbtJtLC3QHLoVoYVG
5C3X5MzIWqtI/egxE5UqS9hSvAk7j82mCEEtL/uW5nN+CF9rd/XST0xWLGqY3qHhppWtiLDJwcVq
8miCRWRtlpJpKBRJw0Lpgvp3R+mCkPwRjTLnQ27uzCYlcD3G57myLM+zwgrQyjTMaXV/a4L5QCcb
ihdX8432BrH8rVWD/ntsP7ydUegmK88zoLWkj/iGYkHZNYGHvSOdQGATOeLvpl75echQPSARbhg2
uqLuzX11FvfecsDarJrMtr1/NFLRMTMYgYQvxlGcKX+LPb4Wk75J94CMabxC1fyLUjHIkLCWvpf8
R8bzubiyH7KfGF++10OzjUXdoKhkrhgz4ymj4hR2Z3aoWqW6YUQJCPaiehb9AExxOv9Jv0OFB/Il
d4O/CHjyeBuX+9lfhqb2XD0miJUbpQqJfyw+CnkhjbAIWOhy+Yw3EGg2kztWrcKvovyPG/i2BYok
ZTWZ5WVK1nbMJOhDPRNf3Lwhb3s63L8jHctNUJbdk2Mm858JjO1/7u07ioCNXLjZfywlW+cfyYO9
FIu1CDNp/ZUNUmWJglGh34gnLuE5c6pqQp+0kZcDWf5Mxb166TzKGL9niutz0uiZoPJ/TCUGZQGB
1/PqDn86lqlOVhh6zjlSQOMXVsyJ3Jz/t055gdSxNffAcciMOwLC7wm+PncCyIFDEue0+8zyUlxw
IE7kg4fzaUGt8bNCnHMmjidyMtSyo7LnGN9infpjIQTybny6t7O6EdKTSkfZDZnFkcXvOoqAVb3E
R5kzbwBQqYR2/CV/zAH58QTq6BY4WJTHLhzyTl0OR3YTVrPpw77kdcclcvWC+hL6V1aSLViw/Sp0
ngGWqL+aSkNl+Rskuzl7PHTa44mxv65dez/SXCYnvK8Y3brvSzzr55vbSDX5KCSCde7zrIgnBZAh
zAStNFu1iA7bl5QmH/1j+LL+5bU0zw5hyWyQIxp5fDHZR6u1IyvIjWeBGGKOmjIXmEJMAUOhI1vE
P+da6vPqDDow50+yvi4Nuc8eeU+bwBZQZVzy6XeJfU34LWrJiDNqUMRcvT6vbTENfo5qcieIuHpL
3YK2jtlFIRQau3sDiyPekCwWWoqH9fUZfFjpmI8n/C+nC8XZznfOFpmWpCdY/lAHiHlbyvhNNhZ8
iqNDk0lIkYIvCkvFWRRjxzOU80qLKXXf4Kh8A7cVWf2jP6LaapvszQ4/0OzFWa7kyH6plM0HdSKw
Yxdx1IldqchhmX1T9WNmCIV11GJDxw+8HT7/tsSjT1lM9QZIb4I/OJ+7q/Bvm4cnRl7TWb/70+XZ
KTN6n4TA6wZf0DnrpPM0YAqOEyZlIVpt2XAf0Bhwpr+0zrJuDm2L8RfYCREZSkikFmZOPrRkTWJq
Vt9nl3MPmyeae5pQFPYmpKwdzbnyp089/VNyh7rrSqHyVnGGMLD/Q9+Yq1fvJwRQSDs7UFa4cHN/
WA8W3RJALQggCrTLAeAVY3d0k/efT5VxGlgJwGbsuOE+PfxHkh+TTyEOC+ElL1RO3T0RgKpsq6mk
C4bBtp32wmPiG4+EN8LrWWjpRA3HjqQT8cqLC6UCb1q8kEfbDZKUX7n/o7dm9EfNqtZ8xpVMoRjj
k/I+CIiGeg82LpbWZPWXPwy4xl6DYSDCs/0Iht8gHXWeHp+j3mP8lyw/iGPw0F0VQt86w+vlFwot
84XeTTwab6F4TglxkQ1fMXhYP4hfXXn1kBPrDLe1dSpKFAVd5UvZBKF50/ULgnq5K7hqCo6OArVj
6aaUI3w2LiuKPZPJNiRtqOuDyIgyLNO6SK0LxPGXohfawZP6mGnZ/JjuTPCFvDqIxh5Nf5OP1sPa
wbN63JNmJK00Q+92d0gbTmpQjrz9kUlWTNGqVsaoagnW0zOEKue6w3F1AIK0iiqGnprEj101mFGl
vHKPA2QK6KiPsnK6WertwkbgbgNIlWjnhMfm9dhyPkjNo2p2b2Ab7lxgygaHMeOj9Iuf9f+Sj1YB
QXC9LllCl7AmoLZC2DFKqPCeRi5a6lwucd9pV0jrhcd0ERYDTLA3i2m0oDXpJcMk4Qo8t1nlKKCi
HNJiapCe5I1JuIajSAV26085OeD0Ka7cRC4fRahsEyueXgyr518p4JSxkYIBOfCYBE5xDViLvDtC
d+JgBl2IABAroYmi746McsvdTQ/oil2rnAEUPJF88hewWPyBicMo/lO8Sd+2rLg+CTubfUJVL+vl
epWhKmxbo/gBmp49AuKeCdTIYCQj0VDJ8mpEzFDTpAF95Sr6ih8q+FmDOmCAQdY50DfYWYcVS5Jx
D4DJI1LTb+8YSWFXlio+EJ9TYXe6763K7lbdklkrH5XcDmqTDbXpVzXyRhCYzbiYcZ3FNFYIqFPA
l0uNMBnHYWIQQKC5FH8sSj6UHdytvydo8V75gL/oCGjPKWMLwdzgxsP2yIcpM3ZKFdFVVhKJXkfF
8LUa/GgfX0M/bBwQsDZ5uqLZtsQj1VyWl7kcKntXhyLngFCLB7QqQwPzY3tXDE0zuVhI9nuMD/kE
SAovjFH18dcz4O97Sa19f8YDq8f+pJ4H9jeOtZYfhY1ozWu/Dt1DvmyGEFe7LWoesy/3nz8KpVvE
ZBd3z/CyByvDYOFlHWmt19suDAOKcpZaLQSGMBAAZGOXrZYLerwWyqfRG8b0/zy9pUTFvW0pBv6q
MqVTZO6KjXfI4VcoF8fiv1/e5TjwVaCq1dkOrzykHIXw9lNnJt1tIMVnQUu285LPuFpweYXjg2rV
nVG1M3xLZ+qSQzof66/SqY+9PQx1/i1Slkqq62EyaG3J3Klz2qLI/vQXR1lWSRn8pV7NW/kiDGTk
vrUTxXjipryZO/6UXHbbgH8N41FA6C7eq3dBoUgzZHqheCXjei1g+6Ryb4QsETB20DFcEhrmQQ4l
qdZJ89c55Wx9IscdEF2kQFyGPWBu/ZPNGIOAa/fpKUb88cjmSPZt335zEjomVA9Y23Jyvq+TLGEB
tIVf1KDDJ971MRC5dzKSeR+uYxox74AVRYGiyLXfpqTrK4DK6fZQKOq73KLIv7ncZtELq7XnFuIv
NkO41JH9ZHXPrgURO55v7mTKmXXvW78NU2i6e8x7rXVm1eK/rkhFwcwUPcQRltXmBSzTj+wbfdOH
ykSU+o+9EMqI+WwtgGOgx+TbRFpcgwmF7AHh/OxbQFaOwrWipv+iIHUeJjxjwdiVxdqpDoBP3eiv
VlnO4F3u6I9cMaPD9MpwmpILjWZvIKCwfivRGhz2TPHfyaIDDjV1PowEDyP7WH/YPRlRSNqNzlc5
0NNYVYhb/E73T47dakuZx+MUHk28HINHKh3aW1qKES5FUTsnuErdVFPuiHl5BvVrNumizGuido9M
TMrZjdEpTzHMzHd0aPqXcKLNIRemK3U/xw5NVeuW453QeZ42QqlvCoTNIW2Osu9eMgrUCsScTlQy
F4+iPAlNpBdPO9kNZVK0OqrnNApWT8Y54r9u6SSCyW2oLIa8SVI6h01l7iYwghmrAa/bN5EG4z9Z
RqycEEmnGck/oB+r7CDpTAg1DUzsZKhD/Bo7P/BOadSgDL1cr2zX7M2o7xLndZh1zSmuwnoV/KZu
SUsFXW9mxeLCZkemeePhsoErpwTaBS/W1C1I5hGwVNHI16dJkSt6Uii7rjiAlcxj155xa+Yyhg9A
WICrwTNmui/bnxsXxsMfUsGTc0j/icvEHdB8XskTo7BLFJ6i0SNBgZZKCzUO7uMIZ5W5vtAZz6f+
Xyu+L4NiWSobbYLivH/kKQXtV8S11Gn4E21Mp1kRkFca2gqhknZOPhkaRao4bqDcZO69iL6e2iXw
dBDA/GPV/kj4NU9+id/S7o9akXSe6+Viskf1Jw7YK80sv20KCSwj7FC+gUlA7/NltJmLrVV52NpG
DT/pmTZem0Hc5ybAfysKkdWNt+6SQ4fb6uDn5Yaq75/xCbXPVeETWxUzkx7SscBfw2vaNAri10iR
rS29+U1pbdYWHkgX5tFOlVBCaIN/msnnV45gyjzu2eWFvpsHVb9YXjuMP4l8DfTx6D+jZmr+5tav
IJmw/QlOArCz/Q4ZLcmD6att8bA8xLOMgJ6rt5IT9Z1tzTRy78Z69+Zfjtl/Q/aV6YQKnEMBllN1
ojIi3L9MqZGoTeejHAdO+eGLtpn4dDtoQ0ADfr3TBOA9K8E1B+mBWNHO1tgWz/gZNAlNB4FHtU9j
u4US3niKQhBQcXu9m1p9EB2uGQpGd67RyOsPh4Kwes05ilYDUPH00i53iJHTpmPkM1cRmSEDn73F
db+QhUf6v2k+iL/fZxs8KyNZ42QU+VTInSVqzlyndzbHvqHzD4zqkReb0mLtbkFIKSZCPnh+Og9W
237Yoi4lblik2nxdgX9JsyYrWqy+hbEcusk2H1H74SgP81noDiPmgLh4jKZ7rOp3dw7WSOOS3d7K
/kRDd/ZfhlYf+U5rSRBypfpyKVgfgPmKOPS6OYG13xF++cYhco2ELz1y/duqrIIwBZAX6V9QnPJg
6N7LkVVcGuN9xewgRNyxMYD00fk/w8+zHCztkr0egowJCfq0L3jvb4gGaWWBbVGFZWd6A/rWxrRk
ZVcnKhs5fNBBJQbevYGraDZB928eJQFbcFvVB/OpG1Q3lqaMWQhNh7jzGHVib59riLDoW9MIGZAX
/3re+gvQ56reuSqpq/Ip2ZhycwQK1IfbAlNKXwko/qOI4h23kK+Wut6rCyXlFlPoqTqFSdkkWqiq
JnGk85YKuiptzaIFJC+vAgxEFaOjYE+uPnhC5U2Suty1AVWXVpKDmN5p+xqXv+sDdU5NmKrdbkQU
UKmwKjK+U/yVIU82Y3z309dzlNrnv6uEt1iHSjWj+gfddfZ2xMDwzyOAKySmWCRYAv3OwpT5nTU4
AN1uKs8TbyZtMaveQFD24rY0Pbvx+Ot5TwDULyJRa57mkUYVbNsO5fFNB4FXs0DoivzyMSz/oDYh
m49rymMnVu7dYvRNK1U9KOD1hkvXqcYUhlh2uEUeVchY3Mv5w5neRf+bqhuukxwn67DOUW9F/0m2
vD04HFcI+aoC4J8vjRR0k0Ijz3dNenq8dio3ltiy2KmCCz+4RU38crpVmUFbVU3FI3LyxRDtR1PP
pq6URFy1SJ+jZk9zX8iaRt9GEHAtJXPjvlwthrbSHBguf0ZZZCvaPhikeYXdNRrjAGV4epH55nV3
bwh/uBR5qOkwhx0gyaFOBrfwRYB728uNt6HViUa/JP8r3EHnzWDlRm0lxbXlZM2dfEjgxDFqOc7r
BJH3jxW6nj/CiteTykK2e29lxG/MRO3Xg5hTR4cM+Km9DiVu7LxfnGZikuoPNUA9MMBRCKGzz1YN
cJq2CMpG0p69VCcVr/NUvk3qo+r2MzVzi0MFGnE+6rR5Bu27pkUY+8XyuIqx7KY+zlF+oKLpC0h0
xt86QyKQ3m/fe5UT//bt1100Di/MhFQqxPvwNRgpNHJNUuG/2tEP4rz5mBMA6hPSgTXNCFqFD22s
kN+OYqjK43drEcuJTaMhF/2e7Efo6bfGzzqy2546EpD27byR63Z6OSFks8KsDFA+2dGN2OrmmzE1
E6tmnJ1nNxMiE9OHGvy/WFg3zWSrTDFuC61L8e6mGbyR5gTvFNk1ELUW5RZt1dttlQS/H4CKGaq0
kNC4aPZjxEAZdKu5HNscOLAtGXwVeZLb4BNRKm7rhwq5KqLSTsL9QrfF8g0mVih1VaOiVxmwNLoN
Hx69kBmhH4KbgXhD0zecqYe1IQR7gP1b+EJbVfrBGL1BSQA82VDKCfAIvVvRov/AahARItoQ0wzc
JvrLAwY4Gru9NEc6ROK1/zqN0aDpZyJeUiVUrdNteJo6tY7pyt7eyLlvZ/UUq+U84LjSI2kqBsrk
sMw2meZ9XRdGUgfN63Q7R/0YZuYKrdHjPsJBodAPM/MGkLdV3e4WhCtzjQvm4dID8beMCrabdxlp
0nkTzxnAp0LcryWojT2zvP8N7yASJtWV2i6bHA0w7qfRdDNlPOtVIX8WOhI40bHEC7atSkS66ojQ
dHf2I61mFcR/o9h1d1gVrZv0EQkWSXBdAGkWYXnZTWjMdSV5KLA2g2IDhoxXOfNr7GmTGAq8EYUZ
bN9IRL3kLzQfLsejueQhi7Kz9RHrxRRLYcn5eXyqsZM9tAGk9SwpsBezSQYCWKcoMNWSHFcgHWQm
qegvBUYzkX8a6SuL9dN3eY/9GhYlg5RqYTLkqdZMAVB0M9xHiEPJ2kHdWGzhSAy4qmJ5NSQGDuzI
lYoyWStaoga9O115VA//NGjIj3z93scaDxpd2JEvsQpnyigwUgDPwBXHnga6Tqa0StnLoBBG2i24
tuRsexyG7iFjotp44N9JAxclRx1u4mmgpsMABbNdz/MIo+xDS2fYPU83Hq5WCoYFAhfsE8G05VWo
3MMhtqm0+kaHyx8u+9wt76c/fZHAPSMnemjZ1kAAsRcEal4/yUEdbK0Lu8mcA7c0fHx8LC5f3Sa9
xhUCZv3diT8fppdM6Ef6qtR3Zw7dPr5rfYYztUxuEhwKV9CSEhueWeEhOCsTdBo+2NMvG4WPQiCx
XS7Gg0v6NUOvMEgDQUleTzAtpepO8vHyu3S11tsSRu1sWQTYKXpQe5qoAQqgygOGi/+zcYWI1RKW
rW/QPYeRt3+7JD1S9GI6/vW8/D34cDYCVORkLx/40ILpc6znXneAqFuNI+6OVIpqt8KaDh7mcHxl
Film0Qu36bUyaawLPL4fDz/UJ+UhJDiVnj2xI02Hc+SmcFu/FKp8dmRRVKw5ctGhgraQlD8jWTXv
0l2gJHwN7/xVY1eh614qUWzcifCOPeebHGG+21Z679RiyezYvsuylq7GX1qEargzpct9582l40yi
BbG8xR3F013+cxPTUnvbxULCPpUUMPZx3QLEz+GJduMhQdn1EyYMdECjtCo+A6VPT2RFEXCdQiCp
KIEr2j/cVYQ1CHW8uooG2tzLr64MTR3lNvCUFR0c0bxKQnZvi/yzgsGVb5PrlbeHGwyP7XRUlq51
zAJ0JM0ZBMzZOhxIHfDCF3xh3v119/VfNS/E1E/KpMYnWhj2j6GEiYSTJVj597umzbV4UWCcHJox
8Dnv4mnwpPMsu7aO6Smx5U0YpAGPENkUhU9rmMQOvAWlUddUP1h9eoJlH2lXkuBq35k/vI8Z9VGq
u8rqznncjGJTOopJawOHP3YX6PT1J9VIXPqZS8VTvgPKeJrX5HpEDyoULHjk9Vg+08xYgdPswUql
sCP5ySAy5BNn9CSstlX0hyNS8ANcOhTXSR72RI4vEZ3eRUKXba7XuzB8NJY20XC3ehN2llNCMUd8
Wy6I9m5nXq2uIxzq4mu6vlER3I1BUReqr4cx6ALtRJwKmUhAHcNGrYV5fiNSfDuZPikdWy5tJiGw
Ri0tAre+e86GmO3kcwu6CJam8JsZfs30zzXiCy1+Pp6w6PTHQt3GXUh7iSGd6NbkI9HPfXsHlFCm
d3eLCf88BKxmHGKj3kHJXbuEIs+dQsrE6DOil8ALS7df977ysXh9w5ovfmVGht5qfkINQRxLLm7i
Ilo1Sik9t6fDS0Ko5MYx0shHGe6sothMJq3jmKdHknKR1KKfnirLTLE3Ql0pWmkwY04L6Mk57eCc
qMx7BaVfbnP/XYLn0ur1j5LUp3wK+T6CZI+7ATZQNrbilPbhX5SVp4PGd/gX9XgZ/11lWZy6Jrjc
OtIJC8g9TJM/4N3IKWH+frMoMxWuaXgDNjoMD0AvqdRtP9QsfOeg5g1c2Z8YNfhzDVy73BSAE0/5
vZ+eMBXGJHnRcOzXk99u6EXmuMOa2v6w8kmk1GNjX/1WMgOL+XqdHmR7iTH6WZ4q1I5+5aIAUaom
0yreX6acfJrCeqmeIUctVLXRNvVHdplmft8Ro3NMr1Qp+FaZBgyibOATEEJtqofeYwDfmcCy3Zxf
EVrIV+XWt7J75xYisqGBLNWuDszuALmtogwG7fUvibXhJJ0A9ZRHJgTtszg0078Z9GzZrjWx9fQS
SP5f8MC6x5jGPhVkHBcrYO19uydxN6P32H3pKsjBF/YcqpFoKf0LajJ5gqKfV1SkZWozWP+8WpIT
k73QlpzVsi3c0vGGj8rAweiXbl305f8GbZt7PGSpDHNHZz6YW6ztFy1iFCX7jAkFCKDTMOmyr28S
g4V32bz7GKF/aXFiVNyDeXDVrr/fzSRJpGqWGgdGY4UDUyF1jSFaBeXqT1pn6k17OCt9lzUFnBwk
2l7ztzcrWYCtFnb6+OCaoQtGgQQjCBY9GIiPfTIpNqu2R73jMA61iQtvGlOasfQehQb8Lgk8wXLN
g/15PipQj9bdWuyBabd9aWGKmi6sCYHBMnJQn05avxkOilBC0hrbm3kCSyy0mUAPcXdAlw/MqpAf
3x8NTqzIkn9X1N6diq6t6rwXn+p5o008sV6ngerzHCN/l8gh1OJdEgRtVnhXQsyckMWK/DERArOD
vgTS6CW5cNkgN3TwMPpRYMbrHFvtVbOJUbjVUSBr7/GpUrMKvcZa6Y0zGCfzog3a2SkOd3xfM+uU
C62dGu4qD4qdGLw1KrcHTBcdtLLw6q0O5rBFJl0slYA8M8ufiAcEGkTa704mvUtNqnaYD93q2KmG
4JAIvfLrsHcBDeFBYxKwNJgrE4CwVGyZr74s1GG8Pl1DBM1NkDCVSWlsP4PdSY1B3wNe1BAQvTTN
tnO0V6b3bfqm5U8JK1z9YEXqiIJbcqhR9wyggFrEJdTigxDIPWzFohziuxYNGjJePe18gfuGK41R
9AUt8+Tj6MyKk32wnjSRHREOX10tm6rWVrRIOZQJ09xEugXDqsTOAq6slZyAJNT+g7FZbYdX3a+7
/mO+jxSWcxwt0SQZA2G4kOIWEAA0zdxCLi5UFGYYOdkUBAfGMWRN+dwiJgLVp1pYoRvERnyu77LA
/t5/eIQTGZD7csMy/ijgrTETUj7QX0TrAGwIDZhCdoJ8/rHY6lczIH/vvha5eYtSy2UZhVihQKYE
rCXNoq9e4uWkxGqFB1UmMCQ1fkJbYv26vr4JxIBBlxz5YmoImH3eVZplqlAkipVcYqVAU9qmuAdQ
6CO2TVULbCwUtPU86x3flZwAlc73D/jd2WPrO786hyIXGcoecceWfLLy2Zp/XG4DIHACFty5iv+6
+dCW+sRvc1B5VMDPQ71d6ADRFkwfbAbUJaU4XAh1ufrYM7RFJKJ9oJxeO4Btz5pFXZjr9iLUSxdL
jtaBRgXclegU1llRaH2pUzPiRpjrPlBL49fBLGWnLdXcOSitE3NVk3T79xokQBr9L0PXGD+0Pm2P
2QRMQyM4u9hAqGj5ki2NcUNh/w45XE6Z/xJxKy1nNHCA2rJFlEL68FwuYxnM53JTiFg5g0AyDTQY
2vW6EtbsBbsjPa/ydROE3X6Mbce0Mt+zvieSmM5y+IuZeuejefibOD2PayQ5uePRqmJ979zxDt2+
6RmiEVVlQuSg9n4tLA7euRzxtlf71AW1akBfDI0aSqM+Ent0TG78UxDNGUEHs4AkwVtq3cq51D+v
eo3cgEkKDFAdxGQSB4JIqm1Q8JtsOB9quNqwVzbL2ye5S+EOWAeCG2kRyCr8G4ZQ24lnrtwbEySy
K6Oj0O2RzyQQTgOY8XT3WZrvvCu2R2mK3poOxX1KYbXoRlwIf8AvzghR5ADbYZj3wsP2qMxa91go
APjuDtDTTkR2fp32zjWMKyj+VvpcejJTG+1pM3H1RBxDP/1swzN4udTs8WLZRIaIhCpnzAO9H0BJ
xhWOQXefvcr44t9K+Zg673Ok2Aq174/AVfhM51GX4EHr6X1ZdDavIL+xz45OCjNuLZ2KfZ8VxRD8
Ke69k7IPG4+MofIuGfmP+3GU8Q/Vr9ojWNuV42vZHA9XruNkhc4f0Q60liW/wuVx2X2NJ2mJfm+f
dKSveIUvx1r2K5yGHLJaLiqO2pxSrc8hxDLTBMj4oi7JZEgTlnBKVuzAMAkHItqNE3yuPK15hWzk
Jx6TVUH04qL4VeRenf9u/oakkh5II0fW1VNgvZNLWH4FXLeHxPvSPisxXUaH7kemWD3cQlrv2o34
iMNfBzhJdXYoaJrlWwOwkXesaJRSj71o7aYGNThIzYqQYvRTCbLu7D3bepYSiPcZh4swNjZLx/46
xjcUs0ZdSUtZnMuXzywa3Pdo//EHrvl3T1C6ukFEE+aQ8YG8mTxej/11o098fJUakZOvyW65u0lY
5yIG1eFna71TNcrGyOII5a6MJMX0LWlZXPglO7ynQC86Lwck8U8lX8miMvE1vVEEtIThdMZcDPLv
eBku77tUhqMzkqGygBjsBnQeOYGkGB0AWPPgk8n9c2rXr7pZ+uM8JRBWL1ZqET6jRBflt6tduptK
yiGhIvxlJRq4cj4g9Q/UE+BTYgm/QMbuysnHKyTUwfGa3X63CF5Rv2CJKllkopEWEkqTrolchMGf
OJfNbflLOsM2RpTr8wblhbiS4VqvDM9ewhWdqo10Vji+dbOjFc2Y8yCLM791cjU/tqgKAwLaXMIs
5P73q0clHp8QH421WTZh9wca6N+m2wBkF3nviE4M0LaRMwXxuiz234CjV2XkciRhl6n06kCOQm9Z
n/eafDKbOgzhFMKoPRN8yAyUks0SRRhDPq0Hp5rz4MiYupM8ofYDGm/47Belg+qUTjd8+CAXp3Bk
11TwGvdnaJBgrkhbuWqEUX+0zvg7MR3D1AS4ATotmep6jfRLjtlMLUAbw6k937IIJC17QQkqlaNn
1ym7ZTZIOTkkuX62QCZagtkMnoPPGuH6waSWD08DeUJIEqRO10pzF29XI+Qb5ae0dkuJAxMmMgGA
48hQ1C77hn2SPkq5WwL4NEhRoqEsoKX4waSz2z9ln4O3CbpW7DcXA/JXLl4DuvyapmJIarPlxjCP
W8ChU6gJ6s29jkXqD7MthrjYhswMwSGv+SW1VSY3iSrhhTwOkWkJT2W2Wi1umGLrlhZbFSG6D827
0SenuXVvCPRzsryrPsAfErI1QUew9uiUtNb1BiQzQVegH1aLLzFjFEaQRoT3XaYtC0sD5IcntHeR
cWYx2Ogj0wphoTXgbJYAJ3nEtIJeFMyidMVhkLUcZY+uWRcKQr1UFX6DIMlnLOHh0oejRe6Wxo5L
MP15LsRGIs4rJvDXJ4JlhsfAzYTOKDdlpfUUNAorNILmQNXx/KpNKcsIHC7mF+r5dGtUFcAXQ0js
tZLk9zJyeuc9dmNX7/7C2/U2cf1nEbgEmq7gnKYXBxh9Nl6zeXP244GT4LoACzOEBo3vxdZtWVjP
NoGG32aOdCSg0McJEt0qvQ0tgnQR3cOcRINqQS3DFgiuS3SkBCjPhD2vuXSHCYjpqwXxlVrFhNHU
l+iuqMtAvxqgiu2zrFsiIQWQH/d6kSxHqoi2KuX4jqQqLPprYsvdxvVae2pWKKJhTfvyTk6YNxcO
mvgfnPMGw3vpMT7v0i0+drCxr7ThlYvrfKAqCT5ITgWE68KipPrAfY7ssjbLgpyJtWgJh8iuFCJ9
nDBrZdSxwCFSw9ZgclXX+BD96/9ZVhGTGVSD7GzQkPAtToGi5QWh+N9wh3DOqdJNM2QTCN0XA1/l
ekXwDkLXsfrt7y3xRZueMG03ITLz9pIO69NPQAdFoczajOgpcAQq3k6yx/LcHVF53QfXSY1gHDvl
B365AvWTDIw09FDKNVVrnEfDmaz7wp4833/NWN7MvBcQNavcBAngi8llg8qS+L9YYn3669bLvg2b
fCp7tpw/tJYVXxE87teyTX+VilqQG55NcXkVYyJIRB//X8VLPWWmizLNmF3f8Lru7E0T0aiMSLrs
1iCmYQkd/AecnLPnPU/bNNYoy0CKRsDQYqtAIYLmHl5titIUvhLboHRjJ26appU3aknLE+HQDB7p
8PATK5r4Usp8+WW7vsPR2lcmt9Idb7XO6WB7ED09S6ecjo2dR+NGcDrEB4n01F7+tXMoJHw5V0SK
LPZgRwADr1VSP73rAGv++S5YmKPWsBZVKWKfkiAEsztYbe+dKnVng1nn4IqGKYTYAOmcFc/duZIY
q66cIe8Y2XcXmn9+5EndpVhwG12gpxVmRU/DY/qnh6MN02ckF3KVAYAOnqVblGr+WwltyqOCB/4T
Ci8PLvNbn6/CQXT04bIuzoMVrbMSs7ZrNw2PfK9Q7j0sEZTEdvx7E+hHJAk79BKa3zDaV7qLxB/O
TEBt3DSsBPjrsfc5D7TwccijEHZ4uYMa+UeR96lBTg8nk3ZIxZlAcOo/Jmt4gj3Xa7UP06gvupHk
cD7ZoenjBIFR9evcgMpbmS4RCjE1wO1GEAxmwKpRV4UAfPLtOcfVv7zY2cshUCpQrOYHG2SsTvEa
1HUAerV88FRRbK0YRJmV0JrLrxnPfZ7pXdqi7PT4iC0ILifUqOYx6zbunWf8syF0tGPIrU40SQEy
GQtpKK9fN2NiunY56pKMnYpwpWyF12UZnP7nm73FS+4IV0joxn8iLOOPBTdBtoD+g3Q8hoNfJiYV
R2+LIGdIVzAT2O0OW+mhOS6ObZGOHDJrPEI5S6ychMEkt7KasKRMxctNch1g/A0nWizwn2kR4u6J
izA7CjEpT1WP+LngmzHT/IcCcVudFgYVsUsxJ5vW7lo2yer6xtZqxF6oTpVRCILyOfKWit+8votG
NLnwAu0uFdCwL44ZJSbhoumM8qqCzX+JheCMmN0k0tKE5xpRDyCdtmPD0uv43JYPIRTt1QaE/aa1
B1ELAHi8JWNRR8Txd49JqeMGmVSAkHTsK+JavRnuA8ovrVWoTZ9JSfLWHhAyklmximT7wuXZs938
W/53WMaShx4CknIrCSDc38hiylzlRyOQH6MwwhkyCVSxjmj/vmeCcMhDgtgFSOUyRdIRrlFZXCJE
A7kXmJRXTmpqa/038jxkROgxEFWuqDoWD+J3Hh7xQ1Fs5aLPuv8sxiNSzkPtcoG1eQmhpntbuJqe
OQiECTIoVQ6cKWFzfe+qGNz/3HbDPMrJLWJ2vC2n1KlxStRDX5Bqja0GyfG5n4HPD5jsPyJM37Xy
k1TSQod6iHi6K6IJzajXbFB1OGMXWDJIe0/1Pamu6HfC4vP+PlPmdfSXh2ZbYXoRedHrdYZBaG91
qHqxZR22zFQLftj+LXsLuTG+tA7ellSZFLF1LRDnanHjxOoIpI5jgxYkmgUI5PBgy32bj0M2LP9P
fK53ONxI8ai6B7Mn/s9BdIexAMz6hMtmDaQzLa5Wx5VjxLEeFYcAVMfoT7ksZJMXQOsBeoOvw/e3
5Vz2ogA4tYm88spNyGv0mXqi+XkpoMc5jMXIT3n0JrLGiEAE1MEE7Iid6+oOZrlNmvo34+/ljhxi
GzXCdmV4hhOwf4xbxKM3J6ZKA5oSHiDtGAhv+LDSJKr68P1SBPhyDYKTeYC+kFos1WT4qApUC7Vj
NQMf+7cRUpwmXvhmLMdSsb6YHqhm3PoL4BOWDvGVLLgHO5XDclouAee2egwmXnTKHB87MpEGmo8W
9uhHrtSEYODPk/XLpy6aqd9XO4YmKAlVW5a6hRrny8Ibu+Ap9K4HhtZLgSbXcdXWUofSjqlWvD3C
v+cyAOhnrpP6ky7sb7l/jKvHDLtuy0PojYVzeREgxb1lNKBCDXeMVjPmOD90ZIS/g6LDWdzDfXwp
lueKhYfEjifttUNJCHiFWrbfY1GRAwrBE4Xqqh4wfy5RKBv2rnp+DP/wBmaszsYYMwvbGcHNg5Sm
PunWLrHNoqKSPS+DpHeA1zrBXOsvwFVReRo8EX/EBY7XccKyeELNn5UQ8PEE0bRzyzSrC4WnSbG4
ZXhRvJe9Szb30AiDtxnqnmWw/o/7+z1RSc4ZGAP0EqpSPxZn4ksphUJ5imaDoF1KkB2nYrlePWEQ
SWZxMyivYOk/h57s8hJ6NjKLWZ9OCi8e2S75ZgquPhkDSers6bUcPEXNwTZPsTzHephNdyQGyEEi
Us9NZ7HVe6xLsnUCVwZvld2Ok0HgfFtX6s3iXXfniuBDlSbhxT9HkGADk/MYYgB6uJN9zey27UV1
4+sDL22j0JPujeBpUmrOqGaFrfJhuFPRvuwMXBA3zdg+ICJMgS9FSONC2IHcmAbIYkrK85775gBm
TdqfqBzZqJ4wZ3Kom/3x3v8PmuKQ2meCeylWv/fNxr6uLbUeRomr57Ru/BNMnntTQi3Dhc+/IA0C
3g38N2vgofzt0hDcbcfcBT5Hz0GcNSV757uA+gTvfXrzErljoPDP5exkrxDbi9FrMa5Jt+e2m1Qm
6Kx9qMg8Iq+N5NZqDfSG9xrdTD30udFBJcYIziNMRM2d6b4EKKo+0lnOR2o91R0GFZjGtGWdKZ17
S9B9JIwCndLhQFWZZYmukb6ZPeHBC7QpPfuwovKDbKwbrXW4nddvG+ZI9OAPQLVrkPgliiNl/VqA
RWeMD7DIIQ9F8nBncLPFE22FoEH6u2A3uDyoINt8q3kSwC21OyJRqiSom4BHYJf2wmbqkTqCKknJ
7hGJpLbQmKqwLCP5wnEUUa8P5RQK1A814c5umnewW7J8tNS6/WkbXlN5WlIrQrrI+bGhfRNe8Pw0
d0hrMjyPZKNIqwFN+KUWzPSGtUzSRJymFEm6srQq967WWVUTAoYbfMhzlICT83eM+m3BbUmr//Wi
6Uz0HouSReEmv4IawYNo+tvz2M1ZoyRSeyv7e8rDjIRW+C9TG360+7voQT0PNeiD4mvH+zRpX7V8
mr+1ZAESkXXB7+KdEhKLSJO1UbfTuMH8JgKCubKU+b0MQ1H1mRMItD9oMPwamqWoD837ijv5c5fS
10BoyWXjvIpLYg91+bUoqhWrHT01queWS6KUL4ukg3/Oe3qvMZdytudz7ZYF2KNNYHSE65VH95rz
F6IirsPp9VjD33BsNPDCokYyxDBWu0OfX0v9h154GNZ0Y2WDlFWaJlnhDdMeE7Gsw0huga5WGPnO
xun4RPENa9xchQdd9gEbREU/6WYZKfc+WsSSJSqokopblLhC4+EtfBryATdk55728G9cfS5CABI5
xwbXXO3vtwkdtagH4lue7FwvSqEyX0MkfRJvuTspUUJC0YhUXj1XFGMzoBStHumbAhMabMkDLmqT
TfZForY3AL447clhx9xiW1ryoNl+ijWnimtIJr3aJRNflOl4wNWTYi1cvtCTK3s1CIo8QOiOXkqC
v8upJ7C5KHopzQkuDsFPDgTlrawixPvdsLLkhuERAYmDHpT1mk6NBf9pezi71eL99ZR4CNnRJ1Ii
J5iEValzNURFGyKyd2iLhrS00sDzSO/hJWgkOu7lMbivxXcgUTd/mq2W6xbSYpj1uHl1c/ivgPja
iOdzzD6p7Pt9f7LhK8xv9u9D/aYSJzWFxGCoUJcgTjwu2iyqeNrZB8L+O064+YcQb+3SvEfgjLna
0zo+zK7N6D69PZ2lnhiVFLhDAIS8QP/ywY2toL/7eOxxPVJV9JowuDgOOnELC/2VdmGcXP6K4FRu
VVWv4eCQd/xAv3rX/cncxf5yN5C+dW64Pq8jQymfws2vzm5uOMOMcnis2TrNgLury8CJ+2Rekeu2
MIM5xNSeHUsesyusO3CeSL2sVfwHiRnaeyMSZz2KkcZwaB7qEeVgvWlLlB6dip2vSKmqJf9LPp0x
S48wQ5C+//TKYtxeBP6G4EnkAtAGKtoAS4SY47PxzGYwhZFOyMk/fjj3fLjuhzcEKGavAIFkoWna
CdWl7mAfmS6h/7CCJDg7iww6rvTQhPm2uUE1bglLiCh9+R+25+GYkmFd30BVdOPS/rvoQgnrkHfn
dflmBX71NALAbY42mfgLvBLRSVP/FBZlxrAgZaN7abDGenFh0BAezU7WS3IkkDlc3gG4Fr3QLfJV
vATKtn87ysC3M8llffWJ8Zx/s/UfCxzGq99/9MxRH3x8ATBaCQGLy2DYXjGnSjz0uIN4LD/Ml33+
HWdwvdZvLQtG/UTFV94e3pcsaMeHNRpDRD4w6wVebDjy/HlYWB7yj+vleLuU5dpE0S+JnnlUIEZH
VlZ7e3MfBmS2hJMsE4/6G83QiRUP8j5Fgmu/F9EriSEpSeIYTOdyYvgdH+S8+1qtO/vk18o7pp0o
OkETu76pTsjDSi77/ydQsxosJDR+fKIxYCPU8siphMz7JeS7bd6dBcHCviXwwyWJj8iCoTXi4exL
0MHNbr9xroS01fqz3NE4P29idgpgrXdE9y1BTIWf6C68LBVyussQzGCSzsRot+zWusEKXx3Gd9D+
35fL0Qy9WgELX/5tgWOI3ChRj3iqdDtX80g98ceMleL9VmuFi9oidCCA4ltOWq5+Dj4Ri5vJKck4
R2MtaLKYjoUxC/7qv0VqU63E9w6AyfmbJNhH3CrEJJp5/RtLHD5xdzjBQs8hZ/i8d43Lm4ogUeDV
mbII4Z9n7VCR0vH6z3vY1ioZED8c9Z1uBiCHUB4OezPBDQyJJaWIVy1/HPSkgqpOz4WrnZMH5LSw
bAWvU1RDU8l9AnQ60TRfNc9vCya7NWEcDnvJC1GxL7EjnZwquktoNs6Iw0VukiXsxKQJ4YC8i/bO
tKDeht7wXZNjW3tbwLNu/8JIhzf8dj1zyC0P/KtDHEPfsEs/GibUnq5EQGPoRaOS8WOMUq41cY0i
1CFDhzL5NCTN7ZdQxC/BobKSIuUsc/nYrUlp999acS9ziX8/NJ3m6qCWnuAeCcgSHIHSk8PWs8jz
ggvVelk+P6X9YHGQjaKyshRthp8lnuSyxhxXGGzrwMb0hzfNjmiIwgBM3s65VTuTEeGYoR2YLt08
sz3AO83ngcIgtgdqNy58Ie39UUDXWLi0gBNEWnb7+1dNDZLETCD7Ps8OL6/dbGTv/TmptmlJ4ama
hhFnjEfcZ5FIVj3nxYVpf7JiLFI+HQsp/ugoslTlbwfIQbOVTEn42an1ZKPh6Pc4akckjmVQB7I6
aaOb9YwTtXqe7e4zU4pk80SCmLTnRbb+Ic1Qqkwi9RfERbrkCff5yuz/NvdTilrjCMOcz1YUEsM8
/BlOidz7CPmKhuEp5LBwL3DEgG3+5son3GPLFxUxm+dXMqwj4R4jQWrFQ5FHgSjJf1ynG6PAwcvm
zAFUtkVw/bTmZcM1VHHz2wusE9jYs1TTT3pGbtceHLb4orRkUNG18JU0F+b9YhG0f316xM01wWoy
ZMcQwqGWBO+fey5FMfst2Go8UHbzTWOXFc81XCzEe3b4zjCVOwrxSGotLnjvLKs4jApsxMHEZW3v
FYfYO1QF5gDrF/8zMKxvmSrbVY3liWIQTU5iSEZ+UMqPnOLPmQ4LSND+h8yisDJePFUVlITgTPYq
bvlznvy9cZzD6kQ1aQFWtI8xSMxAppvqDeeCYHu6jB1d7Hf1+/F7NH6hSF4Vb4BxIWIclV0nxSqb
OyMLp7o2YgF+04jaf7s3I5oPIFPqBsGmFPEN9ahd37I4YDBGzOXqf7BN1S5BvcQRx6UaH49z0lRN
j0QFLLFUvwLgrscmtiCVw0ptCzcFOZ5/bdqFbDtWnOCqL0oWoDroGjoySVNypD4R5O/3m4NB9CHO
U7QFDUzGY6MLuj6RJp3GPOjx80K/gEBXaxrDtz2flZ7xXmVZF/O7qOo6Tgf6FS6SNftqzt80mawC
9VbJ5mlk3VQy/jcxgizeU5ERSXiX7O4TwEcSJOgGrhVLWG6nHLcZN0cTxoz+gOp2szXRGwAPlkQ8
EMX+sk6u7z+FQJdNFWmU4HwWIJUaupKxnh8l8Czr22b6xV8byf9BhiygBWPk0DG5ZwJTbg+FP0HJ
9ypefrAownd8RqRaPIenvP0CV4bvlBcejiuM8BHKqiMzeKg230KwSjD8C6vXWmXwza4ta2YUN8Da
J+puYRiPo9DTxb7OICfJdq7yzzqRxAu/9AuI8XKZF3dtjpm6BUfn6iUJ5AnszxETc0B2qDpGG5W4
A8Q6FSGHvTW2XGZjErga+ehtIz98+nbGQ8pX7mK8wCTQvDeDOOQeDuwqkulW/iqCzRwySGOMht+D
3nzZqtdfHEPvAqVnUW09ckD2j1LHvY1tWFZsm4FJHc5I62WZoIICzEzi/sU8UZK6qycbQZm6U3E7
xj0xKX/NC9Tw2hrnQWCMcQ/x9Ba6lnZH8GcpLNaQgCnr+rdMkbRXyJM5iFZzoHL9MGGwdSATU9Xt
fXlKplvvxKAZxOt93R2s4ug3PtNWHwQkGYRetgwZZ/M6HcXmUHsR0UKWsW7GsmBS+x+tGF6Q9A2q
BVToeyTfmBZKSLZwonFG0GakEqj+Y3jtxPFjMnC9xjQaquiOr14uf9mDNWmt2UJ5XomA1pKvk0CM
cGlcoL0EKfItwIHmKegJyzZ7zTSLc9jXfU3XFZom6LfNYKHdm/Q63tlcImsX5g11wnlUgstgip4M
bceovB1Z+hDr08Ue5IK7OgMqwgLrdfVWed6rQS/80328lZ4hu5dR4FtYcrTFdu27vkcjvWDGDGtT
eh28XNoeFuOGUOwoKXx6aPZhidLJZYZ1lW/z2LywPiFl0NyBEMLaMe2XVKbqHaoTKM7NETmeUiYl
bZH/yneRP8ubeJpE1LLD+v574fWeO+W5fjomkZxCr5swcSvy6gU2KUFBwJol3YAVfy/UyJkCIlZP
Tu1geTQeiv/slKbZDLpUndvKNS3mEBAO6wdvpcNrGUM/5ys7hmR3+vmnd2Knd0x5PcKwzwhY4WCD
iDkBoMm1u2IWpnklyUM5qcMb0tCcsK1MK2ay8txAFgPn/lN5eErrfsynxEYfO8knb9AiO78hA75B
KjQd/CJ/uTTR7UuCRh4zKnMQJmPyAlY0E3OWuG3QQ8I3scYmxc3uSdQME1KsTX9NrsMV6ancKoLV
6aKSGqHCP5okNA4c89Vw13zGwSeSEq5XlmqKHIySN8aFKyhmtQ4mD9xokvyrXGI9wh0nlsdVIl/t
K9e0H781Sg77P/ITuOvtDRolY8mGEkclPU03olsSU9JVz5UiyrNOnU1tO08EbA8GU5KO+Ga4f8zN
FE08q9rlSd7vgUdlLLFLBCgQAD9Flou/zLPVeOWjWDDYPcz4yhORq1QB1hTV5hLXFi805aRtmfeg
ll/m5Tq7xAazJWBvCz26Z0m8ZixOAFyAZuXYGMIWQdFFm66Ay/niIxNGu776Us5ISYPVFH5rElQy
G3/6QqEuXe8hfNqddVwwdaGHHAW4hKiEU5Y5XJ93gNRuZnUJoFyOgAWIzaxs5J91AR49K0RREitl
RI8amVjld7n/59JXObuQX/UbJhrnJ9c0PyejxMw+7MzQlM0/O46+Q8NKvdXxnkWKBF27oh9dvitf
PPBrMImprAsbFaj+Ef6ibcqmqD+qhoHsHvQ/n1wszyjGpZVd1/0TrtNQAHxZofQyQvTd6VYZv1RI
OEdsjS14G5hglv0oUcHyHRaS6kH8H077/WD+n7+8C6BXEp/sPPVetXCCMeHBu3JaS8Xw0T+e6E9C
goGxWEMbTpKdSFC71NppmShFydoL88GdjOP7Ce75l7R6crVxDRujNUwNcve4sEQuBO8TICUpx/tp
DgYgewQ35q63CUedbMSs1AfK0vwexd5TG7h+XGee1W9Um3c4dalSq614WyXIA9giw6J0jfu1a1FU
jwHoeNRMDo1CigmWQ7azlDC7FTAfZocDxGkpBahbhRTvCHPbhW7nTBMUUh1ubLd8uTOCggi2b8/2
vFAPxmodd5+YSuAO2zdedrtjBR82o2vsZXtN+CN7gUXTZcew8N19QW+Zg5o7ygb6BtS/93uaAJIl
qZWJht1fMyUdohGfcYc5r7UnlOGIok85NQNeTAzKvn0CucggKXEvmv3EF1fbFQB3mEp2oythQyDc
EbMM8Gcow9/clhxx4ud7WHQInBNqksuttNwFvJXW5iIx4Xz+UW5dLdB3kAhWa1z9U2VDklO79N1V
9Hp4CNSnfG/N2Jqn9EkwRYPYPGhoT2ohUvF6XJhBlZtgGIFZzWyZafPxCSF3Sabqd/m+Z4JW0jFp
sWmiCXfkYVuxia0x6smuSuzkKjuGu8NqSch0qjzOLzqJz/vGw6ARrEnELyqdA2WoxRezc84T2hTf
M2zgkNnR0Ynt+5Xtdx2Gkyj6JZxpHz/MzqiE1Rtya9mxKnleUi1tDnISvy3odMulQxE6uA4u2glK
EY75Rxotktzaza9FhagABHqo9l49NEm0trIOOsA+tCOwbT0nbRGPpVv0h5Mispp0y0CuVrz5cCa3
zpA0BAIHVxIRD4fSy6bWGXP9kbDCNcTgmnC82GLvH/carNHBTjBYqAiou+c/2aBF2XMEdurNMVRW
Yxd4xHvTNKKqQEOyzEGBb/ons/7/3wp5DF6w5uUyEW5Mnv85V9vDkPLHZP64ZcXMfaVhrxcmZaJy
3s7WgMfsG2VW9Utk2FioVZr8yAEp3nagqE1+ciM3HI4EyWM6zGXIUt/qSpzNPTewHjwGUGkF5k1f
Nvf0d0PgOxscgxOJgne9iub3zb9IlaWPpUiIE3vsylP2lfLEoU3BqwwWhSrWCEYpNDaBbZoTGCOq
XGO0Ske5PIlqXXFeaHdzxjozhf0o4gxgtmyIw7cOIjCjTMjZjfAhSH1GKRbsUfkAxjsdncZI7FIB
3HkgWFWE+caRVMYunIOgQ/Fdtei9Opm+UZZRw96TE7Xj225PD8q491IN5ZSXPo0V6xgeuAraLiZN
P4OclXj0aB7+RUEVwK9KmUuTkjOGgDzxFL0wUHgz2BaVajWuk2konnSGAGjvrHka2zLwdp4rWCHL
PMrRPQT9PFVcnMuX18uTjv/8wQpjZmIiGkXY7Squxy5qo6EWy+igXZcvCv6EcdP+3Fq69JISkc0b
OQlC9LKrJMB8WjHjPNnbspI1eeZq58/W88sK4ZhvpBQY2oZCWYo9qwtN3Nqxf1A2aNcXHN6aVHMH
cdOS0mOQpwrylF4fe94X2aWlc7rT2GlNt5Oc1P9NQDsaKxgWjDqJvgQyGj4B5u266ZArGRfItbhw
bVJDpTNq7izKyBr5TxowyvOR6Ec6f/bOOIBbQ54u//Idm6a7nkOKxrksYhl4u48iLpeL5r66nGLH
E6rMof9lc3g6tkQRv1inPlmtXmrp5aFd+gn0RfThfkvAnpOHBj6b9WEhTwY1MV3spBRlinMUzNIl
acTTvMEVSIu+h8JuXu27YMw7jlnTVpGq6gb+K0LsRZKc5n+NDqvzwVwhzF3aWUZapgTxMiGbCwxW
x5lyvVZTHpy3YN0x5vTfJD/zR1CLHXA+k/2IBrZunBtBg19bPRUB5CTLwX3Pv2j2oo1ve5RYAnWb
AOFttZiuXS3PSyLsLiVR3F4fA4r+NBnii4QO142UdgahqUdR3tJlu0vEZ3EIjxvIkvq1WFQ44/sN
aKU79hDf8oNdMEHKtM1nnoCghg6m79PogOuR5Krk47U7voUaTHq5q+zlYrbwL239uZSfMGeEkYX7
W4dR/5ahmDRoS83UcAjxnGngSlS00ADIScpOAaQLAO3wo858sbeOuSPo+qTa35maiJGyBZF1NaAt
dpWgScEvMWgODA9p3O6vSsNxrK60KX5EGRPTRBXGW9IKZ2RyzoIjPPXu/WZ9yxLV3PfoIpd4gOAK
x0dNTR3OR4/C7ESxtEBceAbD3Z1q0bcfHnT4MDmgSvunntK8tGVQrOrWZhPQU1ykkjhxoSG0M6Gn
qHNzSt/zFQXaga5MCNud1TI0LJM/S8jjnalkOinHwPv8h9YghDMhyaE6vpsMd9M4NnvmBmy/8Hy3
WCwFjGfk97vcGUBm/TEVcLEjr6fhzL7xDGrCKkz8xm0LQ6Br32dPsV+sTtqCHR9dtREMiy5AaLIm
yvwC8T3D5IHAknagl/I+W0fMz2q1i1gAuXTVPnjCE9ItBytndCsZQB2iUFiePv+HpHRFXpTfsiuv
PD3Rcy10KCYT5jU75XTTPpJO9thZSn25tAG0WXWHUJ6jDfNRZgmGprqm80QFkulk1TVmiC5oHEa7
SjhXqwfqAsKjIkDGbb9DbeJnxQcP98B0+71t4suHqDAKvl+UhhcqSLP1tm5xvvtNiY5WW7jOnT5/
ygxDMCjj1rP3+dvJtK2SvLROhs01wl15p0k9vLKQ4Q8M/2ph5h2YObEopPXChcugZSydybdSMDYO
0zO9lzeHCKfqj3LYLas/C78YG9aGFuRQghXhDtxNx5G8g9SgHBBR5tLmuD3NswNXkV3Ewnl3auX+
6YHipjuhQTdipk+nYIUn/h33Svkh9yKvrnvivzuhAhofWrw1It03QwWjlcE2JLLTyMO38wSECtPx
3f/6A/FpwPME4KZz7U89IA7VEabkNYZKa0sLhF0A9nUTDKmX8nx26VB+HNPHVpj58LAKtqzdbFzB
XE7JAzvqOQt+xrFbfwcB3DfMmgpS4p4LBzx4RoXKTbgDHdm3ZVSioPlVf5nwiJZKDk86LcYDs+c3
Pr0mv1AIu991CGpQliFg65FDiGH7CJPPu6lj6jYFhg/qeNF744Yd8MdvsIm/QXrVX9cP71LW5IOG
ir3hezUXYcPJW6tr0TWhy2fd3RIivrix03t8dhodcv2yXi1GyOE08PTZMThxTAqv9hB+stomgJBW
+MJsJmL8qJrLPcVXCmHV+nHyglhoW0/LUvBPiK2UFmk/Zi4GUPacEAgJYQfMFv4nQuwv0a40qgE7
mukI8hLflRP4Heg4V8JSkHZHhXpmZoPvp/eKkMYfMwlHnwMnk3iafBX7G1dL+IEuxq8O4i+yseOJ
2gEtRqQHe5rwS0+BMHWft5fKqdZE2Jmi3ZZNvyFXctF01319fwrvg7ybDlnOybTjFCl/iFLW9VVA
H2Ar3kT5J6Ar3yAYv2veBVNG3dDTyv/kRIxXPn6XlwpcJTxVLirEehqn34IgS/Tfebukug/PcCgp
XCBoydEEkKkmaJiz+5I+es9DpM4PmHFPKFL6AzjjQRljgVD+0osZFb+8tLD+jV2m23crA6Xk/MUV
RU5o+hhd8qBEvHU3Q6xWaHKz6a+q73Nnk38PuWRRhCOr9QKMP32neMRuSgaO7aRQeM5NqtfDDq89
pSzNLpnw6XTXsM+pj9Jld41vIMwlU8RSOljkRe78h2IaXO/HQ6SkwqtRQyu1suWOJY7EzqT64xE8
1t2jZyu/UaRLePifJ/94LI4VSYK2uEnZ0pfsOmpblbiRi3/cASRo5Lfb2M0rwvWCh5x3FnxVGa5N
pKwKQDyT37s+g7s0ZUH5iyH+Eh2IZcwxpGZDURSmVl+r1qXAg2Mb0XLp5p++QETCEaldimcFSgSU
MS7sBDdWLYRAD2skanEkU8sx607jiRvVq9WoSvwW7YEPIrF8jJ6cse/HhnOMQeBKfkKA/l12SWxB
pd/LPAC5LU9XKtlrgXc+UUwzJYzQhBoAu5IMyHlghvRWigDOl0xWk1B5A/PXuJmHDdRink7Z59jR
m0iq3CzEHTgKDBYdQbfzugQsheB4qD7DZ4qKj54HH14c2uzI0cZL5x5563RtH7pFSBZqS80zSoBl
LdbDIB2QVileac5GU38tO0sRzuAi1PvL5iUGnk+f2PMYVXTcuA3RgoBhikSsQgE7tMYYEylVAQlx
2br/5Fy0Wp1hGApnZUs1n0jdjhXj+9ulAJD82jVOLLMwdU4sHNuBITFD5kabJ8tL1nKTjYLBOtD/
e39R0ZTQbbySGZCY44g3qGdYK9aiajbDF+hukQGjOOBq3h7TPjc5WDFDr36SkmTsSc8eNU1MRMs6
WvQ/kC4bicFJFQuCYjuzuEbvWpR29ea94gSidjhO4/SJHysKT7wvEo2QBThKC5gVSlOReDNXkDiA
i3Uue+yeknQHemkW0ps9u7eTi/Cqh8ZIFZr8goRKOQ1jE+zobXe36BzOYA8PUTbj6GxXa8d94si+
cgOi3064pxixz1V/XqUOsxFLxv/2DhEI5czxpdH4OXfJ9CpXFFico27/9F/PRIneCPgv8fi3auwp
xMnI/WpA1Wx0b0Xlj596AmVvcbf4BLEnFEY677wQxF8IyI/kG8enOr8y76/UUdEGxQ2MoUHSYote
05tmYaq+9rBEff2MhW5RIVK5/fBl0YHMiK2JDchI6r8l8kAujPLaneYCvgNP4Z1riHgORtJs/hKu
QXkhEKwRnBfxwuDsUAc+5CJqKT1HYk05ToH8U8n2+GESqN2eBoR2PsxRNPk7SBo5CljzGrH5gUiF
d+une/gXSQ3rFKtf8spN1sbeuwuMxTFZuH3NnrqHmNoh96I2axQofFptkR/pYGtwMyIMW+TczajQ
FAHPHONirRAOe85JdSL4e8XwUQfKPEZkElGvZerk/PoLubqrLhnBkUwUw6fIi+RaTr/Ml7jEgy0n
CqUT5l188HuJYd0dUaH2tHSuI/PxwBrA1iZQSP6uBj9PR8mz1GWKOulgk3u0ke0B7Rps472JK07M
PLkoWvusIrflqLcqzGtLZIcorxlCL9zhWHaHnEkslruyM9GM44uAeSPAFayhvOjMva2VJvnUD/3u
tj7kc3XZtd9l7G2zmlnPjACi/iYzP6cptCbIll24HMIYM5CF2V/l5ZeAFx399Yu7qpgqNR+qWIEt
hPLVWvpfroufkps3Fj5aMCqsP0psH8Fpv7NPEPNMifsMfLh20KbaaGPBWclO0aszzYuu7QEIzJ2g
keDat1LEWf2o/chdAssY1shTk8AXUJTILwnqdwhWMKdqXfzX6SFPUaqWxgAcM8inRIez7p0AEHvf
LDUq/RsSh9JBn3OvSRwF77MegUArO6ylWGKT+KLiPkLv7ycv/sJ83v8zYvjbqUmm4xaut4JWmtOI
qEKukFHhrSAhMbdQP1Wbq4ZV9eITqNb48rpUgsxpzsEISHGx1Wuo570l1fGs2n05tEX2HkWUglRc
Ex7iTe27pbaDp2VXEoR6cD9ppsZ5LWKgz66lEB/9ZRvbkAhMH1tOU5bVeeHHwvEsplk4ir5UhuBk
o1vrZH6lGeymwBoQ+ZLhJJ7JJx2IOEhUE5/SK3HQ1jzK1neLCFzcySy0XiiWjBsqP8VuIxEaSzeh
srMaU1htP5xIQfubgOH1eMuqC4V0qe/24LmQZbX91FxZi7TXKmV+iBotVz5BWULK2FVFk/grLjxB
8RlrHQgSjmTps0FAm5PH3ykp/zuPSxVQb5TbxfFY4w3aFUhnRk+wFQamQB4fXyk7+okQHuNEIE+O
u25/UGBNmsIyQOJxfQQdwzh7no9A6O7LJSmCe3B1IiUfsQQjHFRnsWuCh5zLMAR/JPRM8ZD8f5Nf
2d/jIDmTHwfZ0LWxN7DLYMNrZg06LftVb5wwW6ybZpL7VqFqwRHEiomLjP8Imd7blcMCv3ucV3z6
/hVxlXWMZm85kcwG6GqlGf5xGdW7+Yoi4+AbtN8URjnMNkFFnlQPvNdC8A+ZpoHs0M5pAB05BWyu
rohJE0VAE4Nzhh9cvDJFpcrhrR4WdjLaThZnNrBJANsBwwb7kPxSjYUtXWwT7hcPbNNQW0t3yWT3
rUh+4dn+owqDCO/hPgLBwdT3OwWsJ3PHawvkqYjEDfJ756RjNBhemv6C8UrfLW+o360/Rfy60ZW9
NX0pJJNLJD/gXbqJu5F5ngz+v3M27NW80fpwajKRw1pLDZh61NkQyFRx+SehS3c0ukAo8iSDaX6k
VZvEQf09uyv00/owKjQ/4g8tj2Cz0awMVxpxv9NSA77i1dSCAYFm3HFu2cGItrWkF+JRabhQljTy
KMlzO5JVvQb9BCfgK+nqA8nl9LaPR8ZkJVNI66tuODMi4m1F+jOVz7NssN5zXwOyTU6IBbh6zjY0
zXdzMCoguPome64XhHEgsyr+q0t5f9Yy6ExMuUDX98pwsks3OhATlHHumqj0cO6oPqLezscTXmLW
JI19gvScY8EsUdrNGzFXOFY6LF145Ls2BPWkGbuhQk0FJb8QV4pltPqKvU5aLDIXA8uB7E49ucjM
GO+h2wRrFSmLkCSCqGko7E9mp6VqHrYQv2keczl16HHjskUYOf6lVF3l7Q85VgeHp+Zl/0HVHLY/
sKT9g6XybheIeikrYU+CE+3HUZthcxB7LCjcYhQ/vP3WoAEe3APw29TeshZLwD6HklkQFGdUploj
eykaaIwSbE6yjUbwSAwv/NP7X7L/0Chcri9yhf5jGwbbfOwGylZrrpDHj0Zyy7Xx92RxaGjl730J
0qA3V3P85WPn352BOInqZwBfr0Y3R1Lq6eeEQHZEOSrXiUcWo1sMlCJKkhzYIoQJc/QV0EI73er4
uBN3u36v4bSdccadBHgSa6hlEQsstBBcmOKgPt/tYMbfnk/wnllxTVHqaS4v3aC975iW6FOk6FCC
QN8kBIG2UZreJ7PNf+EbyHFamBQGSFkSIOel/JdpletozaNo+smBcuBtjts4yE/w2cSCE3FuQ75T
M7ajRc2ko9C6zV64EoBYbbiEVIsOF9Lg9sN9wyu5cYcCaA2g26gzdXCGQRv1iseMmw4b4k2F8KLx
SmcnPLrzI15YkO/fp0D/IVn+8+obbAwmEhnS383magcElYnQ+zsHyg7O0+FZEeSrnSe8gJpOCiRK
Ith4f8DYLYLEcPMKpKFbL71W1JzRwVEWghNPWBQjPMAGtFeTHPztuDQwnhgzM99EewbeWsViiUhK
ZqiyCkkHl7sctD58TaasYMhSBDWBJBeQFYGUPGizRyYWXPrqeMa7i7rd+X8dbJdz23lbbf+2oUzx
mgZkdSEAiA7WF/uVa9iEx6TTVo0cCZ4RZ5HA92b/cr0T/KOi2UriTf1Dx8u/0QlW0Rgc9kV8z04Q
OS08pjVwS4GAcRzcZyNX5kmhEgq/n5grewkdfXhB1semlr5vWoOWPiqlckO/cwUrKY2E4HX6Z3Nf
9qYcYQsjmxvY0PGz3X1hYypqZRUNWOSTZPE+gZSwTPPy820z2AJo0ZP+rUNUpEt4eVnjNJGsCFhA
CoZfCeQaTgQ24WvujagIXW/LOrN5Ioz2JzlsE2KKhhOX7S+mCqFiQCyjIM84PjpSjbMsKETIlQUK
0iwWPuW96ZGv43ju9Kr8ARiZYdRXRRHtMyVm7ySloQu6BfdIyd5UzvUb0OMO2spV1QoUhHs8KnOh
mXzfz5gsdVFRdC/ll9ATDDO9qO2v4wC7fgeQ85OSKdNro/cMGEbNmAh9i547thrypQVubnH4/rN8
TcV1QNeLkIc1zqXa1TtQscRlOH6vQP+ovrYWCo3aVHCwA/ipDSNEWVhDls5BZJG1fIczMIiPq415
OiuYfXdI81lA/6l63+8KfR4LUCWdH7HHOSqbAI9RBCZh2Wd4KprK/JraFNXQm48PFzvhh7qc/HAx
3GrKMcRK1G9dDJySTrge4n5NU1lRejslQy4V8praNDYAk4nxTs+KYmewGGo+T3tX6yWir6XVbQQ9
aaHo+bS98d/vP4O5azhwckcZilebJaTVbJCDhTRdn664nfzkzRPIqldh17KSORO8WRUpNyFrrIwH
ZbjEUoWjhaYLz1P5KWuh6YVOSTQTHmQF7idwVxjD0dBAIDXrF0xgyOujxsX3rqCQWZPeLHxRHE+5
H+nWQYmtBmNrXK0PAaEIynDyp0QYw2TUgGJwU/VUyR++cfMZi2WrYDCzV8mH6MoRkdgt53d4whVI
QqpFr3HMS81vQQn3A06km7oMDsQmEx2wWfI+jSDxzV+zqBPf9+FYGSO+crxrlHp0C7NVhZws5aHT
WjPMw8Yjg+Eu07zOSFj1XvMoC4Jku0aYRK7WpBF9QFFK+NPCtPA45TtwpTf+RzycFuWSSNxDx5Co
Ehb8m9mhikiWWyou/UPoWKOmRdcuT6X4xOrquxFadEst/KqMg/Bp1TBq3Igzb+Ts7SfXLs2BaO52
gfdv9DCJxX6U+dzH52AqXYWO6PRmjmBK3rR2RZghljG7ZGPDolEdp5E+TN6VKCzsJFZt2g3iicKt
k6d7sI4pc87VKCibfkicD2YrrzE2+gJxtyPGyQtZ1ChPXgqyCQtX1YXgaqXhZLIrkNWlgrK9ohxv
F/b0BXgNau5dcpFYrVY/t0ko45VTYgKh2CRKPzd19tdfJdmynWdzJVGGKVUWZInK930dRWzz6BP4
PnHrLNX3eRKHIO/s5HISoLu639NAe9SvozUT5zVIP+GEhvUqhyIV65/7HuCJBALFFEEoIfekWjcG
dHGR6j72E8klUVvDN1YHTtlGuXOJ2bOGL9lofRFgcwIE5W/gFEqxnAQ61fdoOvUOm6dJGDe+q6Vq
5CaIJy8360JildQc/tnh/dDn+V2+mGm/CwiqT644uvplgcD+bS2rJnvJ3WxJP7IQyKf2B+0aOStI
qYanfxyZsJw2ry+1LwWkeLroVT/JFgQdHK+Gjp/vbrhjmiNnxYOdGXDWVqntUstZCtF3WoJFphNW
3zVj+mggHG+yjZuOdd5im7zUObv/ksFBCb42j8pzbKd7hEXXSrDO+rEOyrQNvJOyaB8/rACKprbw
nHzfrV9lTi0hDj7x8AivJdqS7EIfnOEDFrtU/b6dKum/0dqcv7vKtTsUm6Kaj0p65FolJBfTmOOv
2EO5B9W+NdTh4ef/Xkte0kKP9igTUR5kyit0+K8vhUHcO+iLsAHfrB23K87ub+J3DOGwn37jOgwC
/OcRW/e+Ky06UMcob6Mnp5NOlPQ/nDKnryZkegNzOMtriADq2CpgKdtmbaTsoijz1MdPvlFaehxn
cixSOgPBwyf8860uP5Osb5YgfJZc5DYP8JGDik2c9IHlYDVJTHNVwWrZQTIihiMttX1aXFD9jFAd
53yVrLs/KCRvU42r1qVmqdcvq2l02xG0Se/1q9WQ7gCwhEAyeUY8NqwOmDCvytJLARvQciUuUv0l
YM3bWnGjOYKewX544ZT8IfSLqzazV0nEjOWEmLhGlb0TMMDP/X/+/OSgMmE8PcyWH2yTksM8lQCg
x7phncnU1nOMfROWLLx8/d8vJqURKktN6+9NHprQaGyoZaGiWl0PEbdo+CGzsXMvH5Pz7ckVzcVj
i4hyXpHzF71Lx09dAgudAf4j2+FugaIr0s+5pHC12iWf0ai50qOKfetgM8ZidDHt6JUSZ+1/dlq2
OG0G9HAMvd8kjNVUm1AGC5tPrw3Q97B4rZdnOEsPFJedsCgDatsXm3i8im2wu0i97b4a/KN6ExQE
Xb7Cg/WL09dXVlUTgrGvr3t1+2zRfIuJOl9iHs7ONODyFC32/3ow4ZWp/SGLkQF1XNyTjhWd2kXX
upZSVwurPzjb5Co853LfZ0xVr4CLacIlqTCGamSa1aRwG18WKZxVxDeIcprVCHLaVp0MLaf4ExbW
GMbxH8sb3vuZeaUeqaFKOyvMde+ofXXeEUPNvN7w62fatIPxqVxpqiLLzgN6cBjM8S+vs4fkYJwf
szfqq/5DkSD4wA/82ocDRsoYSN7gvy2K/MLZAtGCjYCVlsNyV5/W7tzduhK+egEp0VochMHOTpgD
zmq2zdZivH6UQVI8Ly3tWSJGGKfivIBlpvIx94+yDeociWYb9oK+kTpljOf1RT5U2Nli4TaTogNS
HgTp1bdKkBB1vmfxeEZBnNy//J673gkq8OUj4Sb1HOnxZLMhSOZOhlt87sGvjrHzTaGx8xh7+TPY
cyL51zHvOkA17WCpnvxEuX/Lh7mudkgINa4zgczq8bMrwp6ewVMemzX6tZbEsNEQqkjvlPzCOpqz
S7Jdh7ueBm3Mr5XQe53lAkqlgu603tbDWjQKTMu/UfvoLKXFwVl5FWRKWxvu788auB6g1vG+wxBa
+99kWeU5wYB8QItqRE2E3TV+iIqRg4x7u0Uz1ImuwKL+PWH9Un1QFN/VCPnxvmZfa+iw0428lLYZ
ONeT6Ldt3m1hSk4cMTlV/gSCwxKipC5P0VWYiM1qJtPEdcD0jzlK+eJ5ocfQ3BsSEZAG/m1IsWQo
k0VHU33IBbqxTJwiOzT2v8FgNJHfcg8+MW/guTc2y1lkFZgik9LSvVqjJZycj2a8XX7nIv+3Y4/g
hEcRfbEthwSpoBVjAbAxIYeun4fqMvPOfUR2S4ELmj2x6u6KGXl4H3v+Ts4D+x4DDh0v1cdDoyai
nurqB2UTc+7bJpyAff0VENAjWlBL0WgGUwCqjra0Irs7lRJn9n1bPlNPm52tmUBKXXbWekk6QgBm
Luiqfpd7NNmw2Jzua22Nd7I0crBj3iVvQ7UcXgxg/7kt6bZdNJvro30ZRnnpm1neOHlwDoiTo98T
an33xuZc7ulsdWXegAw4MqBuaV9fts2F9FCWfBdHoZnBc8nWTzLzt5XDBWqNWx9jVaCQc1YQOHtE
dccaL29tXrviWyvW9gv7jFoch2Gy5FqfK3cUsnO6yeJgzOYihGJssjPnS9TetsNb8Z13O7b4BBVD
RrGM+gYzLF/CALl2303WJhCfENH2jnOu1tRZ9tvWedpJvDtz31CqtNskzLpKNShjoORqn2r5HRwU
GLZ4qD/1I6iqWhAlAB7AIeNQgyoHmLBmxQPvTheWyVMoJB001KJwWKMUOoAjoouqD/WctvKmUinF
EKem3OPVlYprY5TwDk8BsWpcPSxteRegmhL2s+Ahka6IGDAt05bgQLX2SS77G7uQlW3+8ubOQSwX
KLLZUgj6O2yS1WmUHHfbqdmqJ7tzFObyQcyUPNpkKao0GhRld381R7iT1jBJba0foCx1kFX2BLgF
QiF5D8mXfR2BP2xRkcnO+s1DnblB1GrbntVsqnuOb8H8/ZGRbsFmejfopDW8d3a7ZtIeDs0PXC9+
58WL7YSszWpqDPnUt6Tb8RDar9VvHuXVG21gFpoa/XLYv5oqPp5+Cqgo6Rm2U1ngTa6ZpSF1REi6
nkrYLU5tVBO75u09LrmnSRWT3SC3y6y146uNWdA/74hpUK3O3u39cQ9/LpPzwvAZnRPZzj5hkoRK
/BLg6X0hd+Tx3Z+62ib8EIkyvAGPj31g+lbyJNUwbOQhwm+E19mjtc7mu0NvMplROx+UCa4Mny7l
pJ5uuRBUd9hXV3JljiTgLesv7Mo7/wB6ObgV/9iFFfYO8V6mmt0MKQSfKMwN7dvp6ByTuD4c4gPC
6S2xQwRNaigXedSWlPy6k0e+tyOmKU2LLLEA/ZQKHU8gW/mEd+ENXdwB/wNrBJkb3pdPxEorllKD
Jt+WLaIFNxs/UH+E8TVPxg8YaIyPVtVzr9OB3OzNGRRTkTRsZpd0FoGBEhClM9KXu9F8jGEy1fDg
HgW9rsfc/RD+U53QErKTxXPlPI59Qz9fiUVc9WAkEyt3sN0tA15o5a5YzhE7pQW2eBWKr3mZdFOO
HEe6P2FOsx72/RxCXspsSjSK+fs29mFnBMAocFdc2Z2x8ypi4CCi5sd3zt9Y7olP3kFxbcM/KCo2
h6voN+h9QXLCyhIfxbFgDhx1Uc18aGdUMkYVP0zjYLCNtlTr+F/+9xzC7EGDv6yw7oEADSWGL1UG
bv8DOg0tYk0ctpirKaiZmcSl3nzFNZaP+K5dQ3I2KNNdBXMF4fNdseDRuhOz10lXXwMR1uI2W6yY
sZunQq4P7gROgmPqoSRlqhWf9hs8DVliKIKIK794i83mQuT5EcprVpDDYYStERKvFTZ2VRiyhqXc
f1Dhp7YM7/VYOZr27MLveUxudF2xybcUUMH53j13N7Wr1mGgvujQz18FOq8JUokuCnEtHtnmIR4K
4/r7svtnCJHuYYQ53Kyc8kAte7VspA41Le1wGV099kGWDRfJGVXfbd64NddRgex0K69ApAODm9s3
Dnw7lJ68s+TTOjKHqeehZBuGxz+tIj1HFFjhIckNI/zTH1r77QAcQrLcIDNImjX8uCiBUOjabd69
/YyvkFIxok6w9oOXr8l3shMMUNLoAOlN6X4fg2iDXXlTh/76QaXMDzWQBVdVPOlAk4vGF+EIWwUW
9Uujf7YPjWz+bvbYTNmK+WTQwRzgfG+hFNSJxraE9LASZE+RK/X7o6j1zq56RvYN+f6EmhKw5d9x
PXQonkAKaHzDhe+RjW1pEuTdMPAQNm6R9PNha65nI/WFweNW1FXIaXg5+RVp6qPHj1hfCNsWsyEU
ZxiHR4YUTn2WTNOzVqHbqPXbGa6FCHtXlZp5vfsNAf5mt4qIHmOugfaP5lurtM/3dzsxEnRHBkz+
XMvskeNorip2AHU9KlA7cVix7CnIswLcFFZ8aoXUTaXHMQXa/tqZmpQgDf74PRY+zENVsKkCfsTR
N32rrJbqOa+uC8GRWct/Hc9iys/8PK58E6wNB5w/EX38BDkAd/ZI0GJrJk3052swZRpFk+nVvsy6
mnCic5ps2lJQ/Op+SR+KXyLZZTdgw2/BSN43hIuwN7gOqkW5LZ5QhdRbEQVUC5Tj1W26v6HVmR/7
ydDi6GCjYK4+2p6hzATVjikOTepyvMTGwMAaUTohIR6ODuxArRXdZafsrkuNGBpM1apG9mBBM4Z4
Vy87n6NluKwTgolbq01I7c/usEIF7MZdk1hQMQm+4EjYVqGeuIJFBxdREOE6b/l9x3gT8QVTkX9W
wFWcanixzamRDOsHK8wapq5C79PQHHZ1tc8bgFY1GWohQNWB54NsBsHQQtaknSYI8xyApPPxTqza
0uFJ0JWUn7fFymoeEXhPaKYzdRYRVlLG2DcnhVRkutCxYN1U2yVhvxPoldcLopa4QrfJccSs7LdX
/23YVFwl2VkAFnZx8UEVDitrgMwWsNUIULOshWEHYIqQ/6rvGChoPQuforZi3NdTAb7HCqcuKvm9
1r6pmi4YWwbK5b8j8mLrZi19ioAZ8EBNqyruPjx28ae79DDS2+GNPFi5TwL1sFH68HKiPfnjVgKl
IlfYXHPzwpnLMwNMPKSXomCTLVw3nCLizLSLWd3DQlFMIxdXj+PBvwJqfagsbTbJmNW+NfPecbJ0
Qryo0H/twfm37GTAEFF44qk2UKkbv/kdWt5AN4CiF5Mjjht+HApK9yDkZ4VY/TGjZFco1WcGwJBV
AkrvVYNYFSyh747ac0DpLYMoW5JwBVu7ME5g6oXqBRThBzV0s7MT8np1/rcMftAlM6PfNHJgnowz
mVKfloAiPDAMAmLJk3njR1RdDldsPbahaBzI2GQjExsIaktdIItjDzlRC29P/fpSL2h2EFfe+AMR
F8DunnQ+5GK4DlbqMV42zBq4E9os1qLMCQ+CueC8ykoH6Q/fyuNRiahN67RELug5biY70WPppLc0
HaJq8jP6dXkbGWaALiIxnp7L3cEEhxXumY3n7TKA8UmXWoqvr5XgQ8HoNcJIFX0gDJezE7Rg0ld1
NS4aPd6sLONeWPCKO2XxXYoZrVkN2xHO6EFY7S7LSHI50lIj9bs4M0sukWohRMlfMzz1ixQld0rX
QazAPCNmiXWh3JrtrSjqWRDVsZSkLug4tYHEo5doBWjVUAElmiaBF+AxM71CbnDPi7ELjFAnzFoG
Af7YJ9jm0OlqpRSLm4ZqWWPAEWF616EWKtycbm/N6qewls9DrRD70Mvdu+1o6gHUByDnkaqsFS82
ieq3nn6Iv9OqzrGt57qjNWUFOcu7mW2m/rd7vS4lKAmUqxMNotvX2ntg01cVKmKOgkG7ymNNelUz
WZkakioGLf9aivWUWVq1tDm33ZIephHTokGRKVw4Vcj7amDN7C01Vyn7U3owF+GtAQkUiBUiJvAd
OjTeGCP7qwaFzX44cavAySeOO8SPBp9gmBevfW/g6OPX9ozonVmwbVuTIeZBvkuwuB/xBm0lAbAh
lt1BsKVXgtE9iAkgbTvnrudRvei4+l7U8ILPT/TTmno/Qim2zw5NVSBBbW6dGOGd4UV+/1diREHX
3IwNPHRk7m8nT8brAEWrvpBkIEZIdP13V8NjDwBKo51582H+FR2kOhgTOemH92uVOLguPV1AepWm
fnKt0TNg8c4IR0r5Y2L8RoLVvgSmPYhr8DG66QNFHIlrbTxOBFrY0Zmvmc8et8pDBErOwYj7q3FN
H5NC3ykw/k0mY60RuviEDTL9knoqMz1iG1RpgPJkmqsK2dgJ2UbhrPyZ9V+nt5sFB8hjc8IITlAq
YmKBunm2mn6jga05jFQ7fOjCFr1FOnTAlbO1rSxcgT4Pump0aOjE8bdYrbWrtOZSEk2IG5lsQwzx
eXOMzsmVsBNaEtjSJaCgUbpD+bxXKRIO0ciLdfTGBzBh9fjObDqQHJSjR4luUDvQAfLMYruECFcs
V7k5tnTxlQeiTHAkWVggc5ZEpCuIcBHWrCX8x8Myt/gbYK8HpgCpfebYA1odP4IacEQUReanfcPP
5bMuG+SROUY7Jx0hMN2X0MBhUXKzuBPZlExi5gJElzSFuE8q7msron4hjvLQn6gxyn93KuGdFR7R
GHSPrwdnBVuYGKvY8rQXCzQhI3YU1sN/v6QT767wypm4CTOw6cf8j3hhudO3v/KT7kUXBL7XAIjC
d63QxzW3nXdMAaePk4wh3xVjlwx/HxsvRfQXu+wR2L5/SzGCz1Gtsk8OuBXn2QjKViQDG+FeyYg6
9++7sSy3qGHigxzj8TxWJVjPv0lZUsLIn9Ra5qnFknOz+wHLTTioqBj5busmSCjysWIlgr6Y1bvM
zKvgOJ5TsKEj2+7XJAJJarR3k9W3/cy3HrMxe+7dNkjEsIJZagMMspMo0zEpKBr3yqoklC2XenE9
cb4XytJtXJ9uaOjjSmVNVn6iyKQF0opAAmNzO9Oz8zDZ+kkJdBa1MWCoVxHODjIrCT/bhhFGHlUw
xDeYKISrznOzF8qGcrwssHk4hgdOiCNI9OafR1BsOvJOC3kb0BoU1VEaRH4bNQwUECc/1KJbhHML
rQ/BafG6UxgBt1FHcDqddY4fplf61X+Z3nd6aqBMdDFkbA14dnjkLcUp4yCGs00THHdpx+9/8gN4
a6r6dx44mDLCEEBqAubFf1XCTVvL81xawne73h9CL8eJSe9AGugehVScO7bKwvbusmJ6Pmuo2BJn
NbxgKNr7/LrJGC4D6hz73ZiNwszpOSQtGrioLXPPfsvqaEaYJACGW9gQBcCpAJ5CDm9Qg/39P18g
4CxQahk5YbUEkxPJGUZAWQSJ0csRFylq5dMCF71EqyPcrFYFTEL/QoJbllZVVKp4K0fCALm0XJif
hCsXdvuPNHUFh+0X1j7CfHCBpTVMryIULNFh5VjLEE41gndhAZB+BE2UeyTgMruff3TDjE+SXDVf
MXm/U0GiEoppMMSbqNX/T+lxJgNpGoHPfbcpOdgR24A8PjXjVSe9l4SDLG/7f4ZnqzsS8sIRsL4O
fR/EYjSneThTGquBBR68q6I8QpsurNirsZrzvJQFtE9SWfZfHjQA2NjDBB6SVvsrjPmWZ0xmtAob
cPo36OUVcq0Dd2+VRS9q8w6lc3xmVBVdmBudV8kci12KvL3fkiNRFLk/2jNizUnzzhTUg1rKw6Mn
OYWvzcE0B5jl8F3Tpq3GKcLcVCAL2wS4R6Y7GdDrFh+XuEIn185WOfLRO0RGKHeg35glUogJHZPV
ED8e3Cpxlu06oV9GgWCxOY7SBk3/7L8ARD2jaERMJS6vBeU/HRbsYf/9qseEG/liPJfXgpdOT/rt
B0BPVJF9sYteWUkfsjxZLzyyPfWpatO8YbJVX6HG+JX4aXQL0y3iZ/P2iC21RRbp20Y0YknKofOy
jpVEB9gVa5he3UyOkrxkndJWMF3pioMrfcntC0xXfoblgHSWH/NKomEKQYjKIPRnkFzsP8O85wA1
CuO/3kD1oR8Z1LrQQIA7kM/Q/CXzESOVvtSIPeNvrN4k3ND1D429YOXDzfPkTiNnRGcVPbhbLWlF
5yyVYXDpaPsC54vxnUvrhULOM/cFkjE98hhTtsg/amnf1I3zOBRKuPZZP5FJb0gTnzIMK+ALYNL0
ypazoLQ6VEAS3i403AZFpw4VSK5XZ3F8wd7GrcxpNtqwvtxJgBXPvaChfodv3Hodxo0htP0zaDxN
ThGVajAtNtaZm8yVjNOgviNcmUAm6u+6a0T1boBoS92W9Mc4AAbTwIsvkf6l6PShPUpdFvyREsL2
qejPHy3KptnFKI8rU4urMqkO95RGptgU04VdaAkjh2UEVrtpiEf5FJ45fKX24pKZ1J1ALIpZVZAA
y050XsVbsybgp1h8sSji5iRARf9hsddrWU2bdUj3YD/v+N5JUb+2rxZMIGBgjtx0M/Zx0rBhXJ9q
cfxS2zQMIb+uaCx5B//Fh1VQg8aETlUVtUooCjEZ6p+2MmNM52Z74tlrBacvW7l4zAD7vaKLGUIK
CSqyHFsjoOhCA0fAeRZyMD3TH8RZ535++8L++t2lrO7aBMM3bShhuxHep8hNaxtRg9HUcAaPE1Ek
1Ym/d/dbBobGj+s6K4LOzTMLvc/bgK/mhK6WgSs+4fMMlWmMkxZZrMpIKqzkrks8tByuI33vB2GV
X67lRKGsf3UJs2Nm7MRlfF+CzPrrNeAmOxhRoXDJ8Hmlx/T7kLTpqiWGx/ee7F8/GxZYhA2+tQiK
JfGykZHc8E6SSqadnF+Cknj+kXA6f27OtY2A4w6v19Wq95ZFwBbruh+tqmjNoEU7lZ/UWS/sSkFa
1uIeu75RvajhgZHSpf+fd1hI9sZ4Po5LllDjTp2zaOjV625nPucXEcWNPP4xNt+5DilDK80Dj4bn
yflBUJgMihvZbfqNgCcDa99Ysg/M1lWXfq46AtNtLh6iiXMo0P6D7XBnuUH6ocdQOcoMnPr47syU
MqOrO3zCebX2kbPXGgawUPQ/BGi2jK2F72LPt2Ynwhdyfwnpnm3Hat6tvEyuMi8HOuY+wKtIGF4o
trsB+rK8CgIyfTnxcdTjC+2YuKTv5wh0J/tr65dQ7Hi1ryONuFDHTu1Oc5qtRlJA5v5fKHjiRbEs
XO61jdsH5iZkunHNoGwViJqPbr7uPKEeW/lMEgoWX9QmlG/dzP3PUKRrN+LZ1m3q4tIMIwAt0NbJ
Mfire/pynB+LfFFs0eOBoUplxRf14UVyORcAgzXtUqBFOrAw73FZgAW0gNqRQDqAyVY9Pn2y/5Im
b2+pFn5msSSH8COt/febyAloUCHmbe2WVoufQBEgpB94oxMUm+0kJXhtn7lZ/hwbuiJjvzV1e5C9
LAv5iZXgz+2bD+axTThVkHlOBd02T2NBBIi8EfuxBIj95yASz798dvNIixYk17NUGdJ4o6mnqBqf
p+pLxHopTvaGHaJxC2RFtC0opHV3yn2saSw+ko1iNe0KgDfFm9ZsjknMJDii4PeYP2mlHASa3nJv
+8yJik9m54ayoxlVRHCy9hRJXI+NvgKY2OxIy4F3/VM0Qyyzchg0ngkV8PZIG8ok+5Oepf4C657z
ZT6Fih8zXFlkq+FNIyo9nyYlipw80gJ7Gw9L2LzS1aQQyzOFxHxhVKG4umJNy4Q7djmgFp39K4U8
e3oPVqwI5/ZRdcDVv1YcB78WthVu8IeYrlI+67TRO/22RmhwxPZ2ylvM6Fq8VQlS/TFw/zKzuX++
BlUKnx7Mr5x+Tun4FkP3uhDWjEgDXlPMHGp84leNbul9cn4DPssgztJx5gvD1XuDve8rnuGaCU9j
iurc9YKPGeu84EKFOjYnag8JZtQ2+eGfmg2VV+VDw2NtOlAWJFLYOp0MbqU9h+3E88nAAwJmKwYh
zz4nCppKG2fgjVhrHZ7a4lIEwVJLrCkcGldb/A3F0ZtyBIeAOtWymIJzkg5a2NzhilGKVTpDnIjY
SVNbO+32wN4d1nfbNc3noSufKPW3y9TfHzHHPxW5uCSZNWAy9jTRVkqOHfuf03qXYY4NTwWEHcXV
Petqk+6cGOLV51xAAqFzaGODBS7Vk8NoE/hZlmBsG/4XkqcIaoiPPdp5hDH1vLEDLJR3SD9YeaLe
BI/03QyH6oX2Si/Hu8nDAaT1SdJIvg17c/0iCSVYjoMWdZt1460fMW2BvB57L9Eeu6echx/ZObhu
GCroNqrTKsg34WXvkv2jekU0uDtm0wDr0THb5q7qEwLVD5MyUiCvXlXM1jrDibfsLrOS+rvjBAGt
yq5wnd2tIDrcwm0v4pbD0kIDhG66IqCkw8s0Xl+IfD3IKNIPgkaSoVOzHBQhgvdkDVzIa6TQY1Fo
eM/k5EjMNC83DqSMa3ZX3UyGZBQbF6qHY0B8Tb5YpuXTJn/2zVoXFinyw4MlygjEa1jCx0d0CiPu
ZwkTERkqUbD4Mp1d5QPN0kda5hAhl2UGwv0woy05JDMvFsTN7PWEH6PHjIMUUKPDkS7MJDCdF4TO
a2CLpByn4tQIH3V6Bk+IKQFKSZvAHb5w4qA4a4HTn1btLOKD8WzeNVPXNmKVHccNTBXp4axeeIJ8
sqipWkAnzncMxheceQWgu+0YRwWJp6Reku1YKTPc0+BiYmaQ2JxCvF26LwELcX2CYLuhhtBakh2D
ur07uSHWjJ9IqIdTqCAE5JqLWxGXNZjyPcUNq1ZXWNHNn3yzPsI42MBxh7w5wQqEHifSb37uzwS2
vRDLeK8FDf6O73RmbQYyNdPQCjggaelcC/WSN7ctywqEdRM0OahTx/Aw4EOt41DDcPHp8kyC2vTg
Rd9WPHHJ4GgSZW6h28SdFChboGAyW38XJb1cO+q0R+lMwcUNCp1/uExEO4jIeC5///wxcckHwMZH
BOhIjwSIBc6ie/TnEaop47qWGpQsfZJrMw56EQI3ntY+js1GbKQ6Ss09c8alQL36arxNtA7jM5Qw
77VVKfYDI8c6drq8Oq94RdeCoYnPyQi+HeKYOpcYIwnHpMWbhPaHlGq/7Kwx3zzkWfxVK+lNfx2J
0QOl7zta4X8rN4ijmwjJDAzFsuPwYpFJW3QmJ39WbDHvUxdzKxccMXqx2kL3cNy1tDdfZ2QTb39U
/cKtXO0198QwIbQOrXfuIaIoCuZnsaGWZ2wJaQK0B1hfq1kd4zyjqL/VXb9AZGgOf9Z4KZVJHwXA
G5vyCfchW9wg0mRnjwZ5KWERfKW31iI+T2FstzHJm3dwBAN4vrS7pEbmYqj/MBDOCtZpQwFji5vD
i+e7j2zuCyKjyRRdhbbFK4+YxYNGnTsPEA0LzyV5Qh0fu/064cL+9jgub/W/bg6dHJHD7qQRXx1U
cVZm+cA5jwNG6i4FFvTn1AF4x2wfNlGAtyjyJmZn3boZj3UGCnUY/jVJ86PqU441fL7uJs8XwmMt
fvK3nHQOElTPbJLDE5S37VFP6rJ373XXnufzat7NCaHk0lAHg6cMVbWOauwxrwcisP8df4ablrM2
HGwyVUvVnj95apuG1XqXHlKDLPyEol0rBCBbcNB0ZVBFPe6UIrCZKr3n3QJEPHiT7nDrY5RiMYnh
tCQhVDhK9oKuGKUgMI8UQZBwtVHBiLf/1+CfGtFOAZPNwRQY8AIWFhELZpEDXj0zmdA+7B4gBfdg
4aOUvHnqlIMTuNfj7G7Pbsmvya52Bq4XuO+w+MMoITcCAu0J9+zMx8y6UpV2bDFI6h4Dv48N1iL4
KQ6uiru6+nNTYPPrwrlRoTVu9egQedjCNYAn73O6W/yEV1dkM0avxWGEsozpwhBOzHEVgdORYHul
vdCrfequiTXT78GRCkb02quLqIsRnc7u8tkABff0SA155Mls+Ozn4T5QIgD7lERypqoWrkNGVLfG
Ac35sIGFm/xRVtpRTrP3js3aLjByRmLGONnWbm5dgz7BYsEPuhj5+kmlnma9ajmigbGlx/aBsjTB
iAO7PTVVrd0tlwPeDXBlrdHQA5cyg7C0ppdc1PimCJ22G0kQ/3ZjjvAYZKOCp0rj33VX3m+A4IGb
4Y/ok3v/iQzCvOdYTE5J8e+gS4tslK6z+xJ2oXBjA2dTGnC3D/Hp87jOSVpivejJ7M2ySn+omcJi
oKtpwqcuDNXbYx4SfCvr72Y5+2+VZl1sCOxRMkINgQnNsQGCS7owJtQ13t+8pyAtiRHBFIN3Q+iP
SL+R00wBNTaLusnKbPXzzkG1HNjRFgrhYUaAa8CU/ILJCgvQG9LGNyZBetNJsbFj51f8LdEGWxoG
2dPToSn1NqMI6YNINK8TBQR5Xh6mNUAfJxScJ3d7UBVjOqB1AqvbQwncAwErgfJq74x5KEiEcvL4
+AZOUPfjtNHo7FPougQnUQPHn/ylz63En3I23Xsp2HaY7Zgf2H6Hlx5hq1SqcP/rqtpy1t560/Pd
evRfSgcuiudTj9SeMNClSLjDnvwMTXb3+88kgW1y/AKbG6oGrb+OOjfrqOmy7gQax+L400p1s7Bx
6FyZkyn+O2t3QFNhKS4XwnBtuSbOFTCKmNJO9xvzW/9Lffrg7d4xM2rT8iCOXrNSgRg69GqXOOpN
Kr9g/gqj+HLGbokrCSekLkS5SQdHZC20mmDfawrZq2tIovpD+d7nNBML7+/DAQ0rKVf79xirCoWj
Q+n2jHQ27T7N7FUcjDLSUsomTIasWYbx9aLXMutJAt+lFW1WxVNiN5yzwYxYhoRTCo7iO9WrKOhC
3iLPXXK3DOuaJNDktfoOSjl6JFF57bGBPl4OfV6kGQYR35Mk8wY58eYTg4Z9GTsE3EBMYuhvOOll
6YDNodSY7DjIi1HUKxiNEHQE40u6tB9B41rM6p3DiSEzQ3eVKjnPY1lHFFQhWEy/yAJhiSCjxn35
nxWeYykJ1gs+QWq2bNG5GI+WZEG0mQL889LbsgtKHp1X/dk/hU8yuIP6xRkjE8P8MPnGAPpcjKft
sAogEkHGPV6oSZJPt/r9Y8fXHS10gcjrfcEUbwA1gTytsBmQOaKJI2OVc5RcPeXdpLK4nOogn/xN
WmxnjEId4PK/II1RD+GFYMT4Ylm+ZtFdr66KoCMGkWVMdk04CTpXdS6dPberAi9Wff3hNKlVjwWP
vmW12phMrRG5es9YMxtd9tScu6J/yrD1mcmVBGenh9j9rwcNKflCQoUSS25EIDfu7fd4dEwlbxjd
UURc2LwBJmcAAIBmcqCmjXIj0DCqdTzy5Cg1KpFqxkvsee2u4gHP/YYcHOSV2pmYstBYHeP5Sg1E
F+AYnLg9p0UnWhW8hTH9xXzEphCzs3yVBqjsRO7pt5BPZGHX1Yxdm/JPGlqbB8DAoFxo3cVnHBwt
NI/wpPq/ZHUUavlSsx3znwPBWUafl8UatKIB2PkeLG78CplDNzwDAJNtj+e0c40jla/eeGX9JjKT
24HY84PgN12FUNrXMmks/UbaTYqAKCE5vvwpf8waBe0Q9ivam/Ktxbeo4ta/WUm9d2UqverfnqwR
YJzIx4DFok7AC9UD2T+3dTbvTf+5wCjk9kIOR7C7c0bigSJ/8fbEbSOedkrfzsEwJSmU2Pa6E0sk
crDQLVUlJgfLouihESKCT6fxzl6BladaOZRolGnX241Tl5MOEG1uYwqa0G+5cmPSoiJeVR/Hlx6r
u2B9BlC+CqoL58wTPK9uxcsraBCMHyqQirlUyA5XM+CwkS0XL7iaQMl7YzFuigyiKs6CbOj8ufDV
YrCfHyVSQN8s2sEBDxiM4+yM7oRHFg/M4SQBm8WUHKCWi+IEe5wiC3lvgBwxeqiShaZbjM2ZagV3
NogPDsT316uyQVDiA/NcgMvYOV4uu22MMCT4VM+e4KvucF7k3Br1UOk0+T39Zyw0FV+tgIL5lM5f
N3Mb0Jt05I9aZArU9HC5iFVQw4tuzzDQfts2KTVTmS3a+cHTd+3fg6OpD8pM+VW/TEr/0ggs3J9E
apIOEe3oWq6UD4irC8LqXm6HtdLzTIda3BgZCt16QFWPildbuykQLSEmGjtwQg3MPq4CpkR6ic38
DROkVUDDYqkeg8fJ6A3Kgh+NBQ5W4n+lIquECr3NzKj3Bjd9b+XZ/aluEYuRRUwnDBwsO8GMwskZ
rObMpZHD4PCLpzLFdQkF0w5/ZyNtCnZp2sxfncFTRkgJEHFlHSxOYEGwKtMdSUwNbYl3HMHNRwEi
4X2hpugHIUeKwTWCXsAXbfNUnsMhU6sgTXe76Ibza5h3UwvTGjvJqPgRcazfNqBvdBGB5+UkYQfn
NCUCRdJ8ndEy4o9+pB4ck0HGAMxLf57UI943o0Dbs0+O7pFO8TA1/VyclNYJvQ+qcfUzwnf6hPsC
b40T7Ap6EgjBkbZxmYZZrTCFb09KgfWLwS5tZ8vlFX2HmzjjinAgNh+zDRfg/YkOskS4xaofWdC7
o292mGA5O6M4OVBQBaOcpqYWfZCsiH/AKZqkzkTJwrFlMFFARnZk53NAVhtjUYbdHviwBzgPlWPx
9Ki/DDTNGFD/YMf27lrEfE66wbw+6ONjAIvSi3JR1SIqzOE8n+K8lPb/pwpriaCkZCg3Nk3kpkty
Qk/QkAe/+Q+qeOPW5KLnfSYX/DAXO3Acc46a3mxD3XMgVxnp0bcNYYfUTNQAmpxnP+AFlBOMfuH3
YbykeWYzjMmvMCZ6cMF2ooubGTCT0530HfFhHln9Da4T/BpDV2rs0FQ0iHC0/RUJZGOoeygKIZdQ
DPDs89/g3ryV0qEIM6GzpBqbIdBR5tA1aXgL8+ByYzYVlfD/OLAK9gBmguyB1lFUHGJG/iVZdVlw
FB3I/QBAp8NW9lGScsNSaawKmfAC9Vjl0vTlcfeSPYX7fs3Hox1ret2NvtnZJn3ScqjMxDlIUxup
tqcfNG3GCXItFBrzEbFc3AuSSKCHMYgUFR4WPso8nSYiPwwAzoGoKpjvxf4EYWJEq7Fn4YifPJGQ
p8/iEaloIqpgmPsrP9VkT+1vIyEF2mKzFD81JTXGPqlj8r2vfNOExNkQVtGrOjJZvYZhBW4cbD53
FEK6plZ416QokFPFFYYYD7q5mxxi3XSDyHiz3zFqf7dMrLorYZaL3S7hoU4Kxc3l4SmGLX1qqxhO
P0DMJG7+pxtpg5V8LvXlVN5tGRKuPz7l6l2Y61Cy1iUx3/a8Gd/QbC3nei2OcbRbHIIDgMoiF2bE
puEdxNdYZXfieLtAAtUILNJ8jYKI81Lqu5Xf6swdEnSPDCsdN5EPZpwDf50KgVq/dRSG3YEIcW5e
ZcfeLbzNa3KRMo84Ca36ZbHSxL4W5RBJ40rTNX9r5zNTVogsZ8F3tpff96E0nON3YkJvk2bBEoHo
CO/a1biLMb01AD4gVuUOUIwCCWqs2PpOSF8YbSxQ1nC+gDo5ytMh/bKsgUQ5X/7s+VAXfrYWquDE
Rk0OZl3EmsAoKw7CKR8tW7iFBTCrt6bagieUKeCRcENI+C/XXffNtC9jOsSdKWUJI6vhnFWAaDNE
2Vab7Fw8bkt5ZgH1G/XRZ+fTiotVMId7M0zXdP0UN1baWR0EFm79PPy6dAnHoIwBNQvuiHHHiQSU
jUG1VvNQ+dO0aVVT+Yg/Rz/VIFPbbEz86hCcQZHInm19rWbPwv06y3Zbfrz9XKweKiir4Vv2DndQ
/sMN4uJyh+1Rrkgf47K2wnpAiZ0eYbaeCgwV35WgqKOM8QA4hH8C9TXIMdm7xJFiAmsZNmDdiBBW
l5DZZGM3RRZne84dWNdtFnAMSxpvq66R/dhMJLy6pQREr/uRuU4lqSGoPY4SemGSh35+obGeaSLl
Tz+QYREv7nF7mo9uzEpYSQjmsm7EuwdH/7ZiqfUKzORDbId1wH6oxJtiI4JzdJLH5JmnSQ+eYsby
djtAbTeJar1a9fIwimyLoaqjwNJ7fgRB2lZUTSDADisU5XaU6Jx3RYrcxk2M//UlIlRmM7fr++wB
fxpugBUcHir5JYG2OL8vLRCWEDrujYaXrVbc06zHpvgWUE3jRWABx+fOm5DgNYiPbNGvWNVQ5peV
Fh/1S7vasVzIlOhGinMBntqf9JpzIYccQ40dCcCXrekzVMBYGH9w9D7o7NDy/Qe+V900gLzx1OVC
TXX815bB4Ol/cbb4iwB1RGqUB9+vgaxknZwCE6Ca/5iH9k6Lz84rlEz5zv9ANABYwCi2oELwzgIx
D0iMrYhBK8S04koDLmifGqfBTPvfBtMZhcVbbdaxfBRUyRMBivU9BxJ3DMM+Ce/ZY8rfdqDGZR7Q
usi9lq63An+1BTVdSp2RA1+2CYPMDtLt27zVASrjMFikgvG3rnsS2pPDt58fiodQo8xffaTcSwf3
WdrRlyBDkw2TIrFaB5JzVkiSeLhpK570UXRdz6/qlRygqnGJ239xNLub4yOXCaOZg8xYm+o0LIb0
gDWz8xtXVynJmzvH3MwCzqDkdFWQZQNfmCvuE936ESmwp75UGVnqSzPJAV6x0t27tf8l8yuIxOx5
6s41MW3k6bQJN3v25Cl0C00wptDTE1r6z43x2Gk11TGPMwAaxmdZwX4iUHOubqyx35wlaNhbfa+k
yuNXq1b9pDelg1mN3ifVB9eYEvnK/WRbWK7D3UhRnL9LyzxW+YVhdFpdwaf9+8SuBK2CB/RqXK/9
r4DgB4ySolSPeJdL3Z9Gy7AU+yFvixcH1egmGB9Tj1CTQjxkCC8jaewDLq2zlmuFCe4gvfizpJnz
uKVWxsloh5sTYbLR2kTC3txkND0SATux8r/Ne13jU85tu5Ict8mg+lFliV9oHQRtOBoUg881jwj1
S2eVsstDGD2CHMWQxVeq6gYl6xl1x+mQF4Qdl6BXaF97eU9nOkb0rxokRsmZ2+BYxIKHRschqvXh
ebrKb6Bi+aVtxqUnO30eAglHxyam9OZl82auJCDSWQq8G1CVbPpD6f3wKRkXpdyiqxUY4bvzGY4B
XvFYgh9yQGhY6tVNCdGflit/ZBDZ+hbmOQzsbWG6WCoxs1tMclGmD6Zv7F9CyCcQVB0VQidHZzCB
V/zWX3V4DtV/jlnqTtcixY4oGYoO3QkCiAw7rGywN3IzVqX8RKu9lHaU4V+gliWqXwsF+M4ONHPs
z9Sy9GQKLTK+MTAneXUOODuMwAfjGSi2eYBsiFvv7f7V/XiSpnE6/JwF9+F7tg+ygMsXcAu6sbvB
mhu7Ll2xovr+idLm9wTp1KIGoxJwJEeRqpZlxIf0LOox1sZssAddlHSSk3bwjBrkBmGXtMNHVez2
u+zErVewC2nOalrJTVLSssIMeJJ8iNoQz65pcViV734c84Fd/ZxXtYLnsWUBCdHvAguXzomerB+f
QkW+juThsotOQRBBkioSF3H2De92zrjERlzuetFaMEnlDCqPl/XeI+9MqJg9Ip/+rvXW8opS9Lh2
eX6RLAPMX5PmTS+qDKwoqGuXSYkds7wD07CWeI2x3RPp2suMtJTCcRdTivPnqr4pduJh2I/oT065
9GrEczBQCX9IqfzWxfVEqiLwVsVrfTaEIAdDS1Lc/dm+M1t2WyPxrHi2QgwM60UREaonLnAHBRMR
wbrIG8+kRFrjlAE6Nvu8Cxx+FSdCKZUNsyDNVKh6o0Jojs0oALBFdJHdgIQVW3HaHhbGTWq3VdfX
eia8Anss1Y531P86gyO8kyuL/iOPoKDUkKhvei9vTpqq2ss2zFpqNdJdPyyfTtZvwqrx/5Bq1rBh
syM1QRGtYDfDloTaRpTNL2eiJJE/LdIadzhYIKZ/dmT25Vp4QA/yG4qfn7ltXbiQKnKg7vrC7nTZ
JAePDJho8xwJmx6rza3iMiAP6VrKYSLH8KnIMBFyBs1JECo9XWW0jd5k7OgqUoANiWiNEWMB1DN1
NOx+7Mp5FtpGydmfxd8eu8Wd3tIvtIaIPLEtzOzTxOOFO0uBzKGHlG7SMZMf2FTKtfBsdidHLZQS
9MAvVC99DILfn4h6voQDUxvffLDa474NpVU0anh6G/lniyZck9unPh2pU0TUyrzkJ9nmxoW9GPbk
wgy6AgTbRM43JkR+r+DSmeg7zMrnNJx26uVYl8F4QIzFnKWKCyx9y0KNoIRz+duPAfDs/Nli19+L
Y12+As8rJtu+tL+VxSvexQOqCLA0iP8bRd1wNroCJ1qvgrALmJz4soyHpqLf9HZ6znSQp7rwUef5
jtrvJzV4ES0OVf0U8i+gE4odOKDWPP/jc8jySjSEgn4YOwK59/tFcn+55GKZngPo5j4sMW6/GSgC
fKCX6ixb6PBTr3RAEUCkrcTGHXgD1JVx3d25xpJBt9/dZaoHJC9GT3omUPv37AE7RL3j/U56ucwO
7xiEhC2RZbUSF+vpoIhTJ1epTHWhbVs3y0gU20mnXvNZuOdwDUbmFmohcEXhujAP//pWW5L2SQdi
SYYdsfKEq0xVc/RxoxOxRcPYZskBJpzdaP7Y7Zy7Bi7qqkkwdKQhQQpbM7dmoydOVB4AgJpx6j4Z
ZJekhIwmFEnbsU4f5dp1GAmH94V647BAswIOer1x5HTv7ugYth2f2qxshjLFFWivUq0cL+A1FE3B
wT2Yktf+aRkJeJVcnXF3EUFlBESI0hqoQfHJESSoqMSbHdCCD/4Yon1nkK2s3ZNh3425NOxQ0163
LGETDbKp3+Ha7kLqmjTCNoS6XjAfebJpAxE48fPTSu0KjXP9Zo8nReoy9OdNHZmMNNp3zefB2cF9
o1i3mqlkXr/6iV8xNf/7VhdLnmbcVwsuKs84yeRgJoQsDTIvwUvfF1vJfyTOOTNCJyDNrpog0F2M
5ZIwCTa9YU6eQ2O5keatvm+oowBHjdKUm3KOV0SOwYumYFyioJxJNqsniawRdc46y8mSbxv2jdui
z0asVNDzooXepGI6cGj+EpGVr38r/NH/OWQAKI4+z4ITp0lanqpgkntGmIIguxcCdc3U0FQCKP9R
GIOEsA+vrDtow8Pbx8D4wM7Y7dD2SMhyCSlb6aN39pZXZYaBA2yj0rB4V5DEZ6KiLM7QdXJwDHro
Xx1pmgxhtcj7KgitZWUMdP1FmlyOmVdWKE38pbhz+NVY1cK/kSH/pAVKc91NtO3Wueep1tzjcr/J
OwO9j3kzJ9DILfUygAGze4idhpbhFrBoLYx+4o0TSeG0LlFjQooQsukg/cQa0UL8fMRwTKrMLqD9
XK61Z60asCa3lCbHzGEr4kN/vgb09NGx4vEw4WpM5akDdYREafQLrzE9/2hmBi8tf0V9XvBlOhXs
itMHqmYJzDKSC4kiVnp8UKilzkbDmPFdQ4AFtu1UqHBNJMgmH8qb65rgfJpimCN5gfd5/MxDLv5R
TEIH6szbR2a6XO6eZRn4Q2NqLv7PyQecY1YxWa0/DbylaaScYUeu5PJHCXjokA6ptkpyMDjXt9pi
7+qmCoiLtqa0EUnUkPtWTUqgFpZnNmIQDDY8RTzNM10Vsppe+ymQBIo3TgdQ7o28jpIh60GpECMd
AuJNsExjTghQqjg0ISHoY1k/irchFBnd05vjTTJgpJFocHK6TE4uSsxoL8nlG6Tn6wxBbu/seRBZ
oTpXuklZH1AV4OTVdCXU8oEYroycb+gwcvZ0rF9fpprakFu+1jicumyi4G+W2GCRkdmjSeVzCyuo
+g0Y712uC3cxilW7Bdp1GZxJDGP3g61pFprMf0/cbWjlouegFlYUl5/pa9UcwLfc7zkTQZUg6NV8
GL8OJKbHyZBLv6Ae4X9gOHA3cMQs1CxDQ9jKreH56RfLbsIu8hjTgPGDRO9uz0525lqw+6C/rT5y
QSV2hIO9Ysv/gAhH5cl/njQDYEVV0PYhyqwCpnRsT2AlFwCgWkUPpB6YI4IVpcXkTE4aRSlcCRcd
IOOLkXbf4WYBxf2xHxeP5IpAiRlMLYra1UTI9Yuuqq1WiMVI62YOeR6Wd+AXAm6a4y3+HPybwf3l
/z+jIjfu6gKjGJXvBdTmB7hFZ5ziVpCMT5a4P4fu+MmwC3HA76+T6jr2VmClvM0Gt43jjvOzSGPA
TqLJRC2Jnufj1//gNia20H+uyGyYvsagQFV7NRKGQ3OG5RCk5P5StB348VMEN2OW/fL08a3zBJGN
tsUBX639kaQKcGGeJzxiGODoOsJJ0Ou7aNW/qgYsor1t1XBwBedB7elVWUrqyd7IRGZxLOy9Q8Fr
08/U2Ho3gystwG2gs6en2+HxUO/36iDLMDZnzvPgj/RVcWo80MugUvOTW3L11p8d2ks0ACzC5eZh
y9fKnD5BoKg6whwHtEclnEDAJ5udhHffduvFqMQXXcrbdSBL5A/2AeCNRHtYcKa8L9jZWvwnQaB6
0u87PAawGQmXjQhnqHcrfABfl9eWkF6fec5D+zhXdOU0axF533B8GyGghsBJUCoIUR1FZgfhUlB5
/FfYAGtYwibvwG/LxtKGAun+vwnG2sPI7NSiEXnH/x7inxZ414/Zjs06dtWYg2SexYr/4kWxXbcj
7Ik+z02IuMVOQbeMZYQ0yccamAhoCzkKKCLhO4e4kchkaEjNCdbinnz2Ta4E19mg2Vqfm2yzLZIv
hB8TGtDt9s+p9D67qVudSatoMNQeC0tnXuy9GCfiv4MMiT2PVO/MqViVOIczen16oO23NvJIb1wd
GXUdPlbyTOeEAqkeQ/WSEk9/wsABVmG1ywtSR1clMUfV/5Aar5QP3rxub3ed/2Axz6b+RYha2qzd
Pd23PpHFkp99EdavOX+RZDiSpePYj4tW0drGWCWWcJiCUtRiUb+N/JtjQy5BUVdXwgQXmXD/JVgP
gwkrELiYJHcvv9Pfywmjjtw1MYtsO9Iwi5vxF5ZCcVdSM+5ttVatBwIDrwNQHRJi+eUu+FLouJQp
eOng9kLy3KzFydn8B242lcDyPbCqzo1mqThDOkdb3mijvkzMl2qdk6y9Xq9DCr1PgOSREqLgbIR5
uLGNaIHWgARiuIXclWjOgHJbkAfeKJH+Q4kZjxTCQ9vQ6ArIWs4oXqGkkG18Vkdx0j4sVSVJxB4H
4VrhUfQo6hEUY2mmTshr6u/0V8OFyrI/YlOg2/I2jWcOxvmeWUam0BoLaaoEbI3LzfcGlQ/IdZ/m
A48nrNsV+y2T4nQYnsD1JHqNb4WDWBlrvx8S94RR6bMZt8BpyeeWyWFuxvrtyJM6V5u1QBfOiIuL
DOKwe7XinwfCd1VmPGEI8QbLmeg41pU5eIAe27EhICi+JL2uGbexghHcSNfYV6p0saQQX6tz6Yef
YX3BCxC14/qdMDI4jEtYbT70c14RsYytOkNXS+Dxc3d5AcphvrIhUJyOllMSNQ2RVwtw4SxTE2I2
6WEekw/Exko6fxZvYdqUm4mu62+d/IDXXFDarYUK9j0l0frdC9XSpuaR/Mls+cZk/R/XJHQCLGyj
U+QlZXyCgi8Mjvuwe4gg+uFD1XbmO4WwZNvHu6DHI37vA+4CKeHkDtUqIR2j4bZDOWCxET5u8zmp
BK93Iwo8nLeWnlGyTpS1UcZasOUajdNrALtx/6L4esuVFDIo+UYEyYHii7+y/r+6gcagQZ+3sJ4F
xdj+CcxQu99E/W//rSsPVa0KHKbP8TBxYGrC6k7mqOk+lM2tDbZs63cMoP1AyxOYvYNDZfCbf1nX
ZRDSHxDsnkI5Ow2Lf/UC/Fcm4qgu/yGX55zYVwfm8TwHvAc338Kp3DLYEB0NLq3yagZMDP0mEica
EwR01GAuE46dCYBm5TEpdvmgfAaNRD5csJDavNFTO/3mEVEemQB4InlS3kkP5CO3+5oG/Ufu4cAh
9xwXsZIBQk/Pg3ltElrYIo/lIyFmjEFcqqvTv6yOQSSFDiE04jULgS1VmS3GhBtxbJ2b8bT6/Rfa
Dlma9eEfxzG2LooXfrfwYYcF/mBvC7xF7g6NqbXOZz9avMuBgZo6dhg7AC2AZU9dCBX75P41emGu
cEfp8ZFd/USgO/Ol7SsyXh34T7rYP8CGeP+bN65yTtbfeyV6B2uP/oQNBLdb9IzCCbrVr1b9LSaQ
tAkRyXXF/6gQRW8K2dpxd33Ws/WH6A2Mzm26ffvhJ3Rb7wjGLYVL2BpF21sB7+Mf4Nb2yW3kvXxP
ypKP48AA5ZznznlJahUde8GwC7s4I1idPpuiT+Iq8oWhvX/gT3rta+eMJMY8C8y1gPXBbQVH97gp
Cwg+8fX3Hy91s4YkP273jF5eG7jSoCH2y4RMfaNIKYKSOaINuc48J6jwat0r9fkWf9ZOftc5B+mS
KIaUmBhYSWA/8+fsFEx8G8j8WAXW6rqinb7O5kIZKsif5JdVitsSOihSmQlN4HhwiPOB65tTC+28
d63roS8YbPoSf8lJgn/7ZycgCb/EbNgPGeqGbW1vA0DSeqR1n7LleHK1arZGipGgxxkf1hw7UVW+
flJ4fiLr1HJ7IcWvcXI945LMNd6I7jdSXk8N2Colm6C9r+Fh2fEtChiZ8dSwUuWlf1qkKTc+tMlc
pWtFT+xJP9+UnJYJ5qCMnbw11JzrSwtXotkyvmjwA/9lud1hoFWtHz5uqIOjMHBqU1hLaEjAGmgU
k85t3UiWjIqwAk+G+lfAoSbADOmQWfDHV5KlHuOqAsxgBPrV0idS1r1L8bWp3YHRs8T1/bpjzome
iFRj0v0LypFB+nkSeW8CJizOW9DlTyUV2GCRiYmKDvEDh/4GPXPinZym/nhWsOl6LwdFnLpImIOC
UGbMQLcVcGfrVMM4tK5Z0mFPFCL7lMkH8vK0/IpAPOWRpmEQLZqk+xHlRF888fCtAqawefrx/sDM
7VxtXoejUyQQdEvOhJKiUBUARUHFu1meT9e84FJk944zVQtrGmoiPMCNRhAbVbkFt9yd+sWXkPfc
AJC8a403nXppCojBUmVD7AZxyhwfafPBId0bb2rSSWgB2UVEkYDbGg4tS0yCPq/GIE1mlblBO0qZ
dLNNHaHOjR9Iro7a5pxb328QAVQ+oUIglvXTqQ38xUKZ7X884n8dymexbCgSll+MXHMZ97v8ZipA
bDQgkV26fI7dy2J5xETxaQNwT2itRGZDwwMiIWJmBnGwpRQ00BLjrLTljFyNeQvdt+R+qd5kAedF
z4en9ZM8Tfnaz92kBYwj1xjgIb6HqGDWF4kihEHCFYi2xNkShQcsf/0HMjorJD7/dU+2HaWG71RM
ohaNg97Y1O2Dqxk9elPB+mByRrAxr18jxAqb1aHrDwWwkznNRzGJap7wZfHdLQ+fXOsaXUKOn5GN
QShZOXa2Hzu01H8Sav55bWsZzbOXqYxky/z4tohB2d2WLMlJ5DIvV4RqFQrqkiNqaeQ8wSubz9WQ
uGV1E6OHWQ+BCe7SlKKzyjZNyWo8zJtC3guOq0CA8Od8PiFcmtgD3Gg5aUv2cIZN5ZzINn9y0M0K
jroxybXLWZvi0fpYyHtmc9Mns9pnXNKCztQnIkR/1MNoLcxu9pGYajD0ZpWrNNFmDxAZOE2vMqdA
mGIDNisHFVWhRmXETRR49Qvab/k4fgESbCz4GYzPos72XyVxaxKsD2sGDA1yk+fSLy6kn7Zz0ozt
KfpQ1biPs2L0lnIlwOoWw2v+4/QfZzRBXG/Xl+OiSgsGl93qzPblnLZKpmybDngkGZIoZpoCL8ft
Sdm8Ut85JebF1gn6ZRsIqkffchs5I1ck6RxAjZRL9SUpoaodrMB8sJxhtUcYF9rKRAUZJraSoSN4
sLsl3+oyuXnuOi6Met0WDQE4CK51C2zyW48KXzU3qu6O+Q22++Ays2sMJrsdXE7/2XT24U9LE0Rj
qYJMyh1pgRCzui4t3+eBOvhZ5nSWyNPN0ZKnJWHVetrlxuEOHvQsQQi6HpQuE3usNlMGsH/mM4v9
scO4LaJ+oTs3cmG+wuYkc51mtRF7h8sTR5RtxpUqNvbCZgK5IzzOfriQGf5+Qh4JbqgkMmjFchPl
uGSCM4OzyPs9PFBmL4hkOgHU3Q3U8MZ7+pn1ieQMCXljkmbeCwP6Cw74EdETk5/O4AfqXLdXbB0w
nDo8Gl6JuHDV2fPd9RiGcXHinsrlWSkHOpw1DwvzHrpGjqto1/u1xDyaJMhF05Lqj78EkP3Gki6q
y+hEaqppobWolEFBhF5dZIfr5ZdXdOOerOe616RJe6CRaeCCjfrrAkFxX/cyj7J/eQaVQpjY004R
JzWb+nJyNqc+fJp6lViwajzamNKoI+MieB/UGt8FxXuC/RkoWw69Xy94iaXI+yHgs0QRxrm/qd6u
kpxlAQdtu/Aafk6Kwa3eEwFGJmlH8q5d4Z1AIkUG8tc3f9Qztdcwudhow8v99/FJY7FPZatbOa+a
ZH5JFHxod3Anz3zvlj6I5DPpy/Bn9+mzG+tSTAYwFvCNQjjAVtshoepIA0Kwl89Zm6p80HTlg1+f
MBNPTvDzNXEvHvcdQn7P9TEAZrz4it9p6gz+A+yKWHQLEke6luw7aAWgBM2DP+BTAKMT82+71m29
4y8tlTmyZF93tJexcTyZyORxHGdVPr1fCJ7qwitBRoRZDWUFADQsnnYmcMd0Jtnwl99MV4drlp2F
lLr2nUa50uhbVB+90MindR2vDGiuk0SVXoAP9VnuFKFTDSpb4BSSrWyaeZ+BxIpSq1ChewoiNN+X
rf45Sl68V0yrr+vvvl+PaYGZNOUZtWQMPcW1j+ZDAeKMRIm2gdRiqV1KAKT06xNEqETelhhJEqqP
8eAWnL4NVJCFYTyI5mpLKWT1sZcPnJfosQbYOCCDKXgpMNtYf1NyELSc1BWwZu9rLleT5r4kOg47
R2dC/+/zBWNvGlfIyOlZXAsoQNJmY/ilBPNVkqetrLtrkbU+cbU7PPoN0GD+2BAQKEM3nbRPKbOJ
k5jaW/5OagRrdrdyjVPvE+nxu6kNWs9d2DtN+7VCLWsKgYbdSeFm/e34g+sNYSqwBjmV9mBrHpQm
mLnI1gcvQ3DaSp3LZy1VTSE1PhVqAORRioFXMGiki0TXBk68EyiZoaHQUELqObap/PjVusGm5JHH
lf8Gm8fX5+/kJOXnAjYDZBIDTKNG8pjFgCmpXugKy0XZl45QC8Dk16f18MSVdQE5tMLLjuOiGwp6
DzXfzA0uOK2WDF7PeFhEdRnSXvQE6EFR5lDojsr+RxzJIozHDPvRgpDIoVaJKUrXSIwcU9etS5O8
QyRKdYeCV2W3QKNwqJeC/bNv6WV+jeaxDxcbJk+uOpBd1bkBjQtnW/kVKZQgDUa+xecJ+2PJYhSx
HdtMz1OLP3V2V1xv+1oSGpISpRPPYfwXWVHqNm69yVFQQY3MSCwSnn/4ec44w1DFCOdIpl0ZlqTt
NKC64mglWuegBYahj4WrJKnljTzGvLWIYBBmuL5+/q0TlB5bWQl3XTxZucg4d9z3GwZ5Mzf2tRvy
ye8gb8eSu0Con05tC21ESitHOS30OZbQp4+X82KH3NjmbjbB1e+p5HS9Y0xVTYtPBf6Ycmd6hX5N
XXRkJdRIgenoSvPwCD22w5EQ77YugKmM7I0RAjqI6KFW4Rq3jBX5+j13Vld3VdgV4JWUiGk6C/uY
/dLErco713+7UjzniogVBEbfNY49rfW9NafDVUIpNs6evdtuCrFszwGgKlTLzGe0k0MZiRtkNP27
w+vs1jWkerWzsufUPRxpooUiU2AYWl9VVq9q8ViKyddO4vKwToCUPDvhGLQSKZ0TAOm+wkUN7t2E
hPDfszIdfH5J0oFPfXoKQwdrI/bOA2X9yQ4IAAOuMMYCLJB//x4hX6k0sude/TWopA5uS9Xdc/zc
F7MHeIq217a85+kv6mUMfg1fAGowi5lxIK5bfRcI9iQMxVgEjI9LenrBgI05yWwQE5rDK6+s+iMR
NP2uLSo06VNjV6lAfKUv3Ah4i4axOLHwfkmGJeJRW7mn1lF3RB8BOlQ47TqcQ9FVPkxR0dRTnS13
uBsLHuLVev0VCYD5xDBx2Z6McGBi3NmoHT2SHeN+sMYHHTzKVGHC99iTFvlMQ20aSJQ8MefWkOqB
x/NLhC0a4avMX/YZskuwudcdMG4eHiBqM6Cp6Pih3Un4UjWAv3iNlgYwkaYFJn3T3tAnAysCrnkx
F7hlbnGxDtsUzEdITrGSPwdiyQHbWgs+dUR3ndtZPj8ZbWr7S8XII9R7Lgr9AILgHVJVGCJG9Agt
xp5xEL7nM9ZsTWqd89gr0rvh+ohHKGxcznopCXGXmPy9kG9ZckGC73Uh0KI5l153PdIHIJz/q4qH
SpNEzxedMToBa1gENDZ0nYaRh52CHztxxKa8bMPK3k+UARa8tEKgj0Hl6K7jiwFjYJRQg+eS7HO5
yfFWgdiM6KF/GdYv9C6GOpjTMTbrhJsprNbstmOmXb2jVfhiB9OYhFBen0hCuDGai1HIFZUoCsVR
fnxQaBg3K7LLo+4wV+dBtHuJV7Zl0qWzZ3aa1iFNyRfpCBX0oG9ROiwuvdpZRr3ZCLaH59Gczsv/
SdSE6iYMgKnhn/55CvLP8TElxHGtuRAmGqbG+qyfHTRVTWUwWR+muYZe9CJ6mFLSvTpgosLi9N4B
BcMTdcZPrMH+0+tI6K3bcttZZFZNXStW47zBKAc8XnrmUukgDveVxl7SVbvG+Nznw+G7dcxMUMp0
flKqmmSeDzWMhXL0hSiQlOtZ/cjz+NABILl+gGkqk6mZXx74a6nsJB+y5jKpM9XVek3DKordzYjG
1+yHr5G0sCZUaHjr5xftUy4t2Eohcef3elwavlxmOeFAnjBaiagrE/4NOSz/R4EhoIz76g+wtbxw
b58yb9HBZFJc/zfluEXSyjcTLSLOycZLirttrwxTry4uNKRseCihV5VojXc+T7cHOA0YdhdnWvRe
FHcgfcslmz0gJBkeYPVK24wcV6Q5losLPB/5OJQIZ1I1eiRv3CyrXkW31x98bECNNwYlVAjs6Eln
jzVmCDQQwSJTq5m9R21HYjIh7xD+CKjXWsjGEUp0PoA3gdnyGaUjssHytIamkH1JhIsndqUzwwU0
OZHsMiSiAZpVdRpRrt23VumNtbb12i1HVj1qQ2YfIB+TJZrCD9pBsMkmn8h72+PsoP+CDD7VH2+O
9/JiYCoBU/QqEWIGCY3MGuZQcNPw5Q/aPsNTpMX3vKQxJNx+loqT92L9C4ulCD4HcbGde4O7rKLU
Y2ACILi9PUzi2ocIpvAmgVb7C+bc30QgrwW3/vCgER8qFSyy5bfmk13SerJ8eaF0hNhz/AAsby52
C9LJYmgd0B2ScIAB9ny7b/1LbOw9fzDfvEOlOxRrDovUiYKE1j4ebqsfVi8osQt8l7zuWC1kwWKt
tj2YsXoyMm2RYMcS6Op5rg3CKkE/ltVOtnQaRhtfQhTPzP88MLoJg9yaxPfpRUbQW2q830fl6bmt
GU62qGlkwoT+FVD21t1gcnWTAkBuGuEtCzb+8EUwV3x7/gNzy0ILraskyc9Ajgb5bQyfd8RiVKor
elsgRhXa4NiTJPf7uYW9luBHQVz1SSiVMl8bRETUATdt96Yxh2vFMsUSVcuEgyymLNaN32oOeH1j
9tUttSSRl0OK+UtW+927h8jJjX2QwbX0BUAM5uKvi2ZzbNHKNtz6OrugKtGJEnk810jgbEdNpEJL
8kt78nZBoPIeTSaEgL0zJRlRt1umErM3zTtaYGfGS9x3r91oijoUoi3TZ5QNITvclLSu6b7Lmdu1
9u/EGBJuwlUmSqGl+I6SiO/PwyOGscum7sTp1AEPM2CmuoCt1PGgBulvtWQLPPqpimw0iyQw4fsa
D3zN/u5mB2uw5HH+3UDVaC5I7i4yCysAOvIF/ynF0yJPSMIcQgT/YVX6td9WwMoaEEHrhjZKtXnw
EI7P7EwQ8YFMiJ7yxvZme7r2ciik51HQYclbn3yx2bc5ZDMwW5dn6msHv7wUoKrEZi+4OXFECWvK
cnUOXxVZSu+3ADa7X8be3p3CcfVyve8S5v2oMsQ74TWNcrmflULFn5RETMb8EVbjOMMOPIUrsJvE
dqfmwR+XdUY+uSNGGUsU/BT9VuZFWAsN8ggDenO9rQQiDCqt5Q/huSNFsyid2MsaRguhNXupI1Sv
ihsBS5gxwYJZKT4S+3TTEma/qck5xw7usJv0jFw8XchqD/V3LDcH58TDaUHl4bcbIajt/U7KmO2R
zZ2pIZx0Fa3rFUHiSqM9cBHjf83pOnHZKcF62xl8Txzp4gcnENkhfmrgooEblgUAVbxomj28Uf4x
qqf7AeAajRjenIWou4KRek2W35C2QKa8wkLR8Fat1honWZv9ky43IF3bNS0YTsR3gPDsOU/vXowM
Occ3m/jLgc5l+M2oh/aGHclDKb2lMi0n61WAkqJD5MyEs/w55TvgAy5rFx811SBZjzQxcJNL9enq
YHMMWT3kODwtu7Pe0Tfm4EU0DJbFqx1HrX/sPkqZ6bPH4fraUyI0JGyeY5aYtZ3qor6414NKzbL2
EYD4ewN573F2jg/4HLUtdwNzuuMTC+Iz131LH1Irzl4qYsc9MDd8ul1pSoRimF430vFIRbn1UGba
54qyEoMltV9yqLkZz1E2LMLf47VORaExvST26Y2LCp4sYkLvALnwy4juH4m8rzYZnEUN62FYwZYv
xPUGs9UoePSmTWWaYYdlyhNTFEh5qfCFv7OQgwa4xeY1pkemwFJetAZ4jKagnZv2T9IXItliy1sx
4HYx3YjiG/VTFkpGgpseBPJhsO4hdZgbBFFwFr2ogc1eLOT1XFbkmhmCeG88StpC+kEtUFMYDfR3
sTdwdyjwd7JPs/5z/y6u77Uns9UddMERvl2SdYeO2qCmgXRxBhoyA2z0XfZZ5+NgrXMxOuuj51H6
3xlY0c/AqlwVbb7F4c/AUhYuFiAJrgFTWHkd+EclnBFBBad32t2F5X4t3sGuhlnAfvTUYpcqdZfa
m6uxZym5XFF1jC6ohtXNxR32mjvjo/fCizf738+DPaFZuAzCQAaoGt+VMnj2Lgz6mVqpwLaAms1z
RMe1DpkcAFqcxLIGUKWiTwcikHjaPb1yBlLsFnloZc2GC4CmCNuqyucAkNkckR/prDsG/Xp5UkjE
AgKARvja2xt4U5xp5ScUh49rdB6WwImTUVpYFNrHyv1B1trJ6G5O4HlnEH85lAgB3Vt6/7Jvm3rk
/OwVL8i/sDupA3FxcC4KYDBVTZwRXIx3xwuot0p5GgqQj3sK3zKdddd9kL9OWh2oxwcio7s7LEUd
igaG1jSSolFWFsanrUgL2VgmAK8moNxv4g8I2BWqRfkupokNx7dCrUGhBvz4WEa0RP/e+OXExdIL
rxy5ZPEi3Pb09YXAYPAMa/R6bv6hQARM8URGjUOFwIWeFjWVUsE8Nx0E8hPQSKpSFc9Vh+E83j6A
E/8DEz+kxjkWXPDyIS75rC0wQVlIOCYzPRwmt5wBbtWh5QwCcraJ9PJyhKOGjrhZ+NulBlK7aecP
Z1F11iu6DravVeWkOIofXqdOPiCKvWc8m/9lvWPUj9E3z1p17eA9DnGdW6JDMhtJhp9OUIVIKkFI
ePp7ok677xenEz541LIlEU2qvHJ1hMo7FIeunUyIvrxdLhpEgn8Ml4stuDLLP6o7/I4CuV6px4fq
W154uw8/YNqE94gZ91TuNkGGjC33axYTPq67yC5nmsnsV3uFv0FsMwrYJCIKDA7CIhc+zOd3WzIE
9aCK5inbrUIHpgFDTs2n5egPnGjrcDhPD8l1Sl1kbPXQg2HLJgujAVJiZYZzLSDThUTLPGIsPhtu
ciR44+mSRvEEhsOhHlQkZJ6mVA4UyiT9QhNlUY5AuTuP6iVUzGuk66nqsuKAW9xATLYrd3MSNu1E
+Ec8duMQ9mayrO0v4coLBFsPnotZPuxwbqb6owH/LnhlVyZ7fszkcpp7HL7ftDfcf52ZKP1YA26W
qaIKWuysXCddPpEmncdrvNglQPZUWU9RSgcN30VRqj3ST59UGd617V8dYKaecE2g/9EqTZcIgoM0
/pFQgdEiMHydf0sGovNlL324hDStZQUIJoSi3olrTZokNYAtMosLFUDfZ58XlaL9WcMXeXpqDc5m
MmdjwIgTEa5t3wgVOInFOHWTj+kTtMMUFAerDSwojlu9BI+nM1lHwZIy/t1mJj01a1vFDNokw4hF
Fdlu/kjL4bHCBbARltxglxcUcbPzvUc+fdOr7KiFc8kuyI7QPs6RGL/W2NKAJQfNfENEha8ZYbmB
Bbe/nucJ1pQ1cJO24u71B2jitozE4v4c+Qs9g+ebGFDoR+IXT5QMdOs9fPELKu2LfAbqEBO/EoMm
0K7H7yBmlze5UTwlLMGJbwUxVDt8QON6B5KKbNgu+jgJLAbvI+ekBMc/z4g5e688l4vCOwUBrsoS
rk3jneg9yNt9s17QdkDfPnNZhmFWfMR0hHOAWzh1YSe6D5EIV5WXyI4XAOJ/FckVbOqoRMlj1vyS
S1GZs9FYgW2fv665geQYsyEXmbmii+t8efyk76t3uyd0CLfRABz7OVf4uuCZ6zbiSkSEfi6Dmchc
j6cOBHuu34z1BqE6/tz48BTK+h0gOZwkAnEtj8aDpZmkciYcoYBqBBZoyjREa/LsfRdErLlMoFaD
chViNlbpjEx/LFlSnuNohr6ASS8OhImY15IkO6iUbmOz5yEj6kF0m57/TYjdurNT0L2f5wn6ed1t
wxR7pexyDtnwH6GZQ5WsXopqFN7sWaVvgFspfqWhVddN1bkvsOJRGFA+xPnTYIjqgE8o/L97pc96
4A/9I/KeeESYWcunyU8vEZtcLwER9Z75WI0kpB7Sk01ePolNoVcD3EKSk4E/ZJp6lVdvvD4PD6jC
8MlqjTHkWfvb+0yPBgdxQEQ+snMse7v5eDRTK3d/Jc/weZyZn3V9cO+bSIk/mIZOqJg21A4UTBQA
UApP5+ghB+2ymfFLzrz4yZxD8y22SqaMYQXkDwhg575RtRSECT5WXWiNFvt/XadA8uuYUAzW4HuL
Sn0t+x2ug5WUiSy/E6/gkRjPxPP4zswCNj7imTuEOXqHyFxCqC0K+FkWiMvWOpBbPxjKBN1R/2zp
qTaMXUcKZyTN4dmEqScFFzREDTVI8u8D4gjL3++A6eAbcY+CIGhzRXL7wYvtquzJUDKNzu/eTQRC
Y0h0qzpzQ7JXw975c9OvNjE4t3nh2/oei723Kaxlo9O4zrgokME9q9lAZTl7p6g8DpR4TPZckupi
cDwx8ATa4Bp5/evjZ8FteVCKpLKFkAXiJ4MWvuieFmibNr6CPsuBH+mq3ssD2tY4+2XnSvrLrcjU
lifDajA3ZjsDS4k77cECJov6HDRAeedpF9C1JorqPHHi2GTM5nlQUTN34YLUjlNmABxUpv1fDlMK
r8SuaSt9gB+BrkdjKTXRtrJKNohYrvyuabVdKmPibG1ehr+Qr/ax6r20Qokh3mZlgl8/yWvPoHqx
uv5LFME97GzI1eUSbPP//XrOJ4CfreL1yK14WTb6BMpaGap3GctZGyY1Sd3a4QBrXxbNrHju6tBS
zKV7/M9q5bqJgXtzdhUeOPNLrGj7Ijs1VV0djYYzi2zutlNQBNXLjjLg4H/H8a5QHPaCHEkDLemQ
m0Q3KuALmsOILGl3sTrUwxIUeFQ9Khf3VB7GKnGDANilKKQXhMDJp40IdUyI212ygn0Nu7GSJKPX
hHWNkJenEm22qbB0cRvGLL53QuypZpZES2Fjwj9ZsiwZUvn7yRJNdXX+t59f6vYWkIobnHQ0cJvQ
pWeif0CC8A1EmpOq2GcULkuoqA5zS49B6hOFE7CKdij6koTihj4XgcYvI4Mzcta/kF89LBxQqlo+
J0bEyvty+UM+GUYh3wJmHvWN/o6Qcl8keHDlySIX/PrERyvn/2x9B9oeRXd5i/wlpH+2I1djdahG
LOSbgYxjvg3tjIo68oOv0pXtjFO1CHsMGnsqnFstqq1r80wyD/O6YsCYFoJCoLuaGMVR/5yM6g8T
ITdouHhUi/7r2Px4PCaUU/BXxmQzPbJAQbaiEkaASIZFMDL29nP2im7Qxs7ww7Wb0Iu7+ksgYZll
jN4D3xcGpyv66QVj+MmFI/++xcd4eTE6YI+scZVVmHyUETCblIynCeEF8wcxhibhb8SojAGjZ8rG
H+twK21si2LhJBYJI0a60HVSlM69L7eniMuBvRAbQK4UKSDO4nLtxyxgO+ClvL7BSbq4rQUT0BaD
H74smqFjX2aHZrubgAtqcEWzhBCq449gjc1qQhzyMg3ALYJxzu7CG2dP2NOIUb9nWJ28/TkPOUcj
NdtnRqCNtw33teK+u2mF+NdiA0B/vCDrFhTWjTW9lJSPansiY81v+aE8QyVJsc5kKhLKIGAGTxRM
ywxNApVQucU3Qa9v7YjJZ681lN5VU1U9ku1kNKvfSoQW4iWobiAkKykFzo0CYqttLQjSw6IfGzvA
iYyzTCBwnSt8DPYQcSxetcvJ9N81ZgCoVYsqtFdA+gUi5iHOU9Ez7yfMp+IwpyjQMrLjXz4zJB9u
FOysE4PPjByfgSbt8w4Q63weQhYw5i9b/Es1WxEaqI1Su29eedvgDgMHypKRAjzgArqixw8vhSbk
i8hzyVL0xhxqKbBfhJCBPsVzpcdAl1Y2tt2xZcZ6VJ/QvGhUPed4IqGrIqJ0GR/3Bks/KItk8LJM
duNp5mYCD7nrn0o+UE9qw6KOgzVRoVaOo6JEDLik1Cc/Th3+B4+e6zvNTP39gyHsYE5A/+CSmrkx
ik8YRMaeDx9tx/XPwA1OD+LppvPWwmJhz1WqZUYXSydnz3V0RRVohMmI3H7ocBgbIGmcRIlCWNZD
nzuLs9Oid2t5KyH5GrPWmnfu/kBwA7ZXgtF721apJaIjRqKruojw4wDEvMPnl5egECsjyXnr8Q48
T2SbCE8GaWeRy6GvDYXYe0GuZuHgNMcu8uIiQUJD6Y4O6uu8etVj/4jMdub24nEeq//C9ohxfy6V
/09owRtNEYlBj3um43d+rtoK1F4SZN6TA0+17f6N5MDfa53gWPUGZQlhYfLuaYLgG2drMdLHf2NA
70rDig4+aAmLItbV+oWpKySB20nyDATO4OJhsQw4XUIvCzU2N2mdJbTTWBBwEJWjNxEe8pc0Q4c4
ooztJ+5Ru8a2xxnjEooW/iRs8LNzExofZQ17yhRdV7GPcZUTUSfAIginUj1mOVHccaE2OcPhJZ08
MtSjgpYOV2BBopinjokJxFeHkda+b5Bu+gcYU+aF2v+vbCSo+9yRTO0nilviTiBH9Ss40Ny51Iuh
kVtVpguzPmGKVVrhOv5CJmSh2dmUrA2qX/xaGIThyqkWet68bybkskbVXr7t2rnlMldCGN+v41mL
BFNqHRA2/l8gGlXeiKbC0jRsSnKeEkRz94MrxiEbEfd4AVWy5X7rt1JXFESSksMdkhBlt/X4/w0F
tFCZoD1AmLEV/+9xOmNXv9COniMm/CCwcFvp7dgAYd1fjcX15/me9taaZZVw+Sd+XMujCm2Gau+r
Mosn5dMgH1nS8DohhXjBPp/SLS0fphmixieiK/QYRfQmUSBiF6R3F/eXsAsNwd3iO9KR3Z8fsUtj
1k8tTdOqSEdPqtadzhdEKOLMheK8DtTSZTR3b12CdESqlhjf1PUTdj17FIf4d6D8q305pe6bQ++5
yehDs/+JS/QAL/vsY0xg/Y0zC+BtNaH0O6CAVLG7iuAeGQwFMtYdZ5pYt//t7f0GT14e4XZte4Jz
HXQ99X6AO/UDaBH2yxSblBwkVQ/4ea51rd1UnShFdbf2H80LjsUM6JvYSc8bNdG9RvvmlrVe7uiP
e6HrhwhwrW/cNbfDShGXO7qeBLqkdNtEVTsCEmQCKxK4AKYdnazTiW1W7AiVkQLD3qrq1LJZ5ERI
PYRXRFwa2K+AOSeuvDLlbUkIU6mlYGB9/ytdR/tFwjFbC+Fu3gZ6KPEuIoVBRhrLUEQOJ42kgWp7
YYeVsgOduSi3thiMXABqGnzbloeLioZt0pi9FNN72BMtOotTMhFGQ8CRYfcCPQRww9V09G9Nhb1j
GG/Aj4O8k4KpjKAFNx2QZ1lnDBpCdvtV6Yxip/jv0ruDafOfTvKRkX8F0+XzD9Yx8Zg8rpE9LViH
7fjRcvv8xXFBSzgU3x1WkKP3WdZei4BBIAFCH9Zf3NzlFM2ldDwRm4B9yblFKc6tgCjNTchpAydq
EHzCAC8dHm2lIVOfoRpd8zA+fhYF1DkDFoXUKFrTsvGPsE7zSY758MGZoM2OyiiOPksES6wR6zeu
gYzTpTmrsAf44qFgmKplbj+b4CpZRJxxWY15i9sgECe+MWRTuyTOGjKYr5xLhPmgVTYJdWgBFIeQ
F1S4kXK7/9Rg7+UyfVvi91HBYr/xUq/g4keNiYU805wtCuu2MZlaVTXBlH6mosZsIiIFSa8DNzU4
gAGztM7McQRfRXP4F3gtBwSGKVtUZG4YcIoLKsw28/IhjvhY3beiXDDbj95ESDhRTqHA8qVTKNgC
w+N1l4CI+uAc9jbwCOKaJEg/krQSSf4lqoZHIwvxEsYjeMvE/rdWSH1KwlKXh8zR7fiMXvCKp1pM
7h4z877wULzn4sAnqKtzYQY851IeVfn13lCeeL/5fZnQPzJ9/zhBcqOd/vytgdPNwMXCIaXRVz+l
IOxidd2JWLspwhgRz/4skhaCvw3Yc08TodrI05TqekhqWteTBH8Hfu9u6sOFv07/C25HM4Zzr4Fy
En6SCvSqUNc/zets0sx+tmGyDEAFsFeCvk8s3iupmHNNdF/jBUXh3aKB4alkhcGccq0SR+rTN4Ym
YnzEDIOLJi9DHC7t6DUeKJ+O0dDadIr9lefgmXcEDSDRrBMEb87OK+7iThoM4L/JVGdOlb+piEqc
BcBPHuuWEqaqGPOQZpdJiv2+mw2DFjYqWbwBZay382q2mdDCR0Cmc4ynQKsT2GjqvnHVKAZfQ8tB
hRaU0dyxAc51z42j0OWMxvZMUKzhNWpT1R746w/TrHQcCCLrTRBZcqkJDBULwCDD1iK7uTJ+r9dx
JKCo2iT4AqGeqRl1hA3n4KrTtY0lNzyENpbUE9CekU3SHk9x9/4whUAkKFbA2Sjhrla8QThbp1dX
ZM/6q+QG3L9S+4V360f1/L2kU2E8YszifsumoifsIHFMed2CxFsS/wLOhJl7rJZTJe4lAdgL7zTR
xqqEjFwi9Zf81pXqfEtUrB0qcmBU0jLqxrRLhsz4ei2rZ0xFJRQdMO8XV4ERjHmpbSp5MmbB1LTv
XFk4P//MbPlBJ/SOuvvWUjfi8sJJ7Ienw/nA8+BrX/4AV4Lo770JBG+iNjvA8+8FMAFXyrVvrys1
pBM69hQyR0pCQl0zOczeXwYJHg5YNy8iflJJsr30i06gLb/1ybCy3uD8MEYPhkm7l44cZUH156um
+YV/KRSPGE+oztQyQNeyXiDmBjT2vskuyHbpZaudS/Vt5x7HVS7Anj82MnhM4rb4cHsnZNYU7w5b
2eJ44tjshm849TuyqcTsGe2NElaXuz5t5f9sxAkI96E+S8vF0VfLftwjvmGJHaYGaxymQceOX+oY
9BUkFVbfOt7pBwLPqaIlvek75cxDq1whRjTsT4cZc7PCcm2RKd/4EtEOZyZ59AcTPJul2oUplj00
TrXdrriwAvXI4IVK4+MblTB2Xo24tYr8bW+/Ncr1m5Y8Ly7OnA2za11k5wCqjhpoJb8VkPUoxXfB
PDalFRThEpcCobmhIUHIA0yhhAfIeNmv1yhtP3iE5mFC2hZkZM3lOz1tjVkaXnYEBu8Zg1Z6+S7g
HI2m4b2Y/VMJa15NAA5udL+zxfgOj2CVYDfyn2HaDZVh7SEwBisBRHrnbbb6mVrN+G4XNKWt3T62
aEJ6Kivo7eXhjJWleNdCM23O1azBxBZn4uwweFrdjKodIfbkdZhIxa//+yhSUymGl6s+//Za9I4Z
Vj2RqMkUtOawYlzJdOw1fmqqHkLxpUIcL00QLewpDKtSBugRG1Y6FEMR5W+uIxU7oB4Vvnm09OhH
R5jiUE6qPnmyS/VI3H0X6qzywKak9jypd7JsoGO9UdlTDqXf26x6TVwNHJ8WfqcGrZooaKjCOaGt
p4eKxjlGDGFCM7HUHusf4Aflm7smFZT4I6Rs04sVvH1lIAm6FgmA90OEnd4mVe1VPQ9c0G2M3sTS
+L191rkM/H4DR63+Ap5bSuaAefLn35jSBvFY/9X+ISt0lDOrgCVlwX9Ue8vT0POTstldEuko/1/I
NHuKO7k1HsqhfSjLAUZmPdH48/zVueLYpgJLpENEGkRnr7mx0s/z+jz2ORO0VOfsxnngxsZByc3r
p82t1WED+tWmFV4RdjaXlfZvD1WGUyKWC71g6cS14tMlixCKm8Ga2U59ueAPR82AvMfjDlA5qUcb
DGNzKqaFPMRnSgCAaziGnljU2LTHLAvz3aHmNzJEuTnIyJOCHWhopRWzq8vTyVKN0arPZsoS7qAx
ATpEg4FlDMCxvbdOY2TP405k7Q7mx9x25be+1eO9bSDGCcdIBfE3qXbG0qIJKvLIGUFdmb7GZCTX
+zrN07yWeS1ehEdG8ItB0S51yWBaIFFXqFcIxo+ztB6efk5odF/0zZ+NOLDBY6H0het6khRpCTh3
mqOHPZiYpqVqryzVSPO23UP+qe/SSqBK5yBiBUkFW9SEvEMTalEBFs8U0afR3w/jRWMMFvQMyRyQ
S9Ja8O8aYcyBdi4wRLh/UH7uHY84ZVxf+5sWxFnvpHWKblE3nIxOjnQOfhPiKKrtnClDOEiDpy0d
oiHzECrrPju8Mc8gNASkz2I99ikVUttkiUPq0ngvUv0mB7D+G9/LRpSi5WktXLGTo46Jwp1ZqTPx
MgZcKr74xNsiDJLSHx6GGYKMsYJfMeaVZcPmF1WDsiAKj2CZzHJwe2feww2svepgmSri8Ckdmqyi
34Z7md2AEoUm08mKL6aOQElnA6mJrc6bfKYnOcXWofX8/XQLJnfiaM6iPT/laydWBoyID+jCdwZw
LiVn5/GltLowwSEUM7F1rRd9gy3WDIdKTFSsNe0oMQ6CQlHNoJUDNzZ+uXuftYnRKwUJVMMRbZlA
yd3+0PV6C/M17qSXTT/8QJFrz85LcqqdQOJnHmL7hylNZa3h8AllET+IIk6GBaxlcD3AFK3Zzqxi
dqPdjyM4XbkoK0PZ/WwFEOlH1O+P4y6krnNyBE68o6SXBm7uj3qrVd/XiPXm1hSLoUJFYKRYygr1
tzz8N5d5ufjCaUkm8w9Oru5+Z9VrQc0ZWt1M/bxj3nRXdNR0Rmw9LNmKh2sEzj4X+cwRF5CAKB6h
fwTJceQPbKdg0UXCG8nKgTTROjQi5ux/DG/MXkIejWdvSYZ2Fq13bwAJ7ZAebBnQMVJ2E86Hr0yt
mPN4jkjMO5r3J/u2PHLvhbLEfu5bicizLQWAWflmWJzd46+BBnU42PYGmDqE7J9F/OYgOrVrxtDt
uoXUyMriU69jju96IzQcwdUiqPfHM/ZEYUdl9J/WkH1XAd7Nzay4s3eIVPgMh+j8LC/Ex432++La
Yihci+13cTbOTAs0tEdhgsWr8o6QFupKt5iQju+xqLnj+7jfTblgj4vWqjWBFke2t1Qxw/cQAqiu
9hNDz8dM9qbcjpUrNxfHPhz+wk/HuLio695TO+eSNdN0v+CvEzIsnlnmRiyPuUrcBGDEs1TJK/8z
RvVs5VV8AT7G40vj/NuTnyGQK5xghlqZJQDHMgiiNC9DSOrWwnICLZVN03mARn/VF0JjAsy/DdkE
RXcMzMLvphenw1STbZ/V4zna1BFqft0DNQQhb3wD5E3hIO/NPhxojDLka7Jhjv/qfCfgIBhbOVgm
Ss0i+7Pvq9MxlXZZ9RhZKQV1pwbfFxiQr/ohfAhp6pjM/hOJIyyiPl3H6KGhnlzCrOjlHtB5e5Aj
5LiekL+Hs/oWMhsFpCZd5F/BCHfXHjdL1UW8ywXEv6S31nyo1xzn0YZDMJXWC7ADyKgOlD/4IGqn
YOkt0UlZR48HafSwa/1xFO+3dLQ/QhRrWicJ4P5OAdkkEsFoS05yGPO5WFXU3/bNTDVPCVSr7D/1
B8eYUSF3/ublBwQ5Cj5WeCHlpsjV4RSfhLYvoYt/qyebZev2QJDo6AbCmDKT9rCo27alEp2ZvIuO
voYOlIK0U3Ox3peFDauOlkqa/oh+ErsPpJDd4+aWdzMX8PEHidl8OvcvQzB+zJmG65fGgTEojKWU
Tvo65lVco4L/eDHSvhMoiboNE1RPFS7jvOEC+iMS7B4GJS2h1fQ6dZ4soLDMhpcR1NgdEFkGuLhZ
6cOHAqiCiUnFolezgEkuapEDbN8Rg6TBM6s6HbHO1rTJ5FeSxi++yG+0kAAyEjZUrlQjYFSl2/1t
TL8XbguMFo0eFDrcryMaVDvs4YtHvqG3Zgj0Fze4x621TyeegHoqt9zlokW660GaOznMrBNBjLxH
lyU/R3zEE3hFTS49uh1SkFpg8huHK5F5PbwOFVXo/zN4DxqxG9P/jQGmntv+1jNzSQpiHvu0TwxD
9qs40jtn1qOx+NTH4YhjtcTE0PX4KD1Tz5UIhYyf3Ib8WHf0Lf5dLDSW6y0xQOt9CIKwr4ApJZVV
T3hoF2ncP7xVuuavYYiCQUkBLUxAi+OfQeI59l4jnlDhQlC/k0s4FHu78mwU4GVyHrzwHDAekClQ
H8wNoDA7Us/+aK08oMc97G5bDSnZKjX9OoC7DHNsWHYckrfrHsn5+0ml697+nX/cs4cZtQ/a+rrH
rNNCKOVjRsDxIQRuzLULWKmvwsCdKla+osMjjhFVIN7JbbzFml53gNVwjF07kMYVCAGH1oNEJHPp
tZfYyuvgAyzXGMXN5Tnd81fR+E3Nd5JwXIN18GbRn0lTsauPsN6+uz4V2PuUenl8miRMhNRiREiN
UThWJfpOkFiDIWBAc11Jc55dq5D3qnHXb7mVdevZGzc7MrLIIOu7tpcSIbZ+/NC54TpwB31yw36k
sVMDZ5+l0qO3qbNAP9RBszKwf8L2K6pU7TF3ntJmFHDMsJ1qLBw+LWP0WSJO4Z1toXy9G8eEgn6v
9DmAkFRbAmrre4Xbus+MMlFPW1sqkgZd9JxndEDwXgRPmFi9HhumXdU7zMMPYFBOLIb7pb0B9bgY
ww7kTZNy1Cp8eHCT9LcZWuJe8AU4+mQbQTkENFeRnFYs/u7MU90TNj2YNpjPVg2A2nCPec+txG1Y
2795HncRWFd2MK5/OZGggH2YIiYjDf5GuwAPdbKctVe01bEAoy53VnpywplROTH81S8mooLZuW3C
Qq/En9w+pBgfYun4SCR57L5iW1wGxTGSKSDuZGX33RiAqCD4+QLGqO30gr+KwEBF7DazyZIfeeuO
cxtg0beFTNvB/PbppcsyDT6xU+t9rFpzR4jBchZ/Tgq6oMmJuMD8S2ERWRFmxkrI2B/TrTwRoRmk
Qbp5GeO5HvuzJAxFz0yEUaQwUYrbqyJuNT+vNE+hFt1Go/ZRoMMouscUuWj0TWf9rfmsFUl5/285
78Q+HPHRK//Pk4rbNaU/kmMxlhr+bo3S1tvJF06UOpgSxotd73VxLztKsduHQZ3j4M56zBIcNIQ4
VtjYaSbN2FZ4Aw8nbx3JslnCGjnKzLfag4yMMvVD4Qa9axJkaUHr0JXZcYFJLDkYTnzTG8Mh07YF
WdvOfzjBZxRTkeHZPWR8/Yypn7DZ0uxfqGaWPsK4J+apnLTp460D8qtD54a8lXzKaO5FTmdqREV5
ForJicAPlCP4wMyDZvZ69N/DMBJIeDKfKq9FC5fMaWI8ZjcT7N6RGBN2vsQqBBazjEHFQLFHTAjE
FTVDKYnrlRALPzT8NSkzkb33EFfjEaJm2mh7pzOPDzoUcJaoGoDmhK5bveF5/slQYWg9XUSihoDN
gTTkT3Xa2o2D7SXPcZwlASQmBzn7Gkfkb+Cl7w+H8QAtDGHSe/8p8N5fArO2vcKoaKu7wbV442Wr
ZuzzQq3TwYHMVwkWTXiv+tOMal46wC9MJvkMQkkeZyqDIB/harcXw49xEQIOFsmMZgWo874k/nOD
n48jVvPPbC+E4sUxoCPiVuHIfBAyWvwNo9MgyET4Lv37zgOaP+GwInR7rScKjHtL1AerhLADYECY
hkjG4LUJaRTzOHvUufCiw5Nf/XusQBG4385cuIyl3uB+0EAb6zao+gC9FVcnRJmNTC3gQ6gnw3EI
rMA/cRcaXpxiA7L20PLrE+N05WTr88JJDH+B784AViTrb7rG2kjGcwVXVzlqshM//JSUJk3K2JA4
CdaQ6GerHjdEKlLwiDKG4EqpQ6vEHFRBuFHfvkYO2Mu6SMrnYhn5vvFeMKoj5eh1kw8fLObfoXjJ
lFojKoJUjPDDQ2fnMJG1Ny1qkactqhrxkVa12Klb4IcEkVQh7a83Wq2M2jUQMx/8enK2Lt3YiObt
g3b5kE7RciJV1Xkxd6PWEuPghq2pHxxJM81NQau1eKjWq1JPivUnqd6bdR8mad3tns7WR4WM/S0F
qNE4vh26+Cwm9HltsL/1rEAt+N/CciMDGbmkZq0J5uXcFeoCt8ULjIbMXkzeJSWBnsAMBvxb5E5q
dL+shf4N+QomU/A+0qGncAmNiozlpv5LjAsygipZUGXn86/Ri3kq/Klx0zPND1JPApP1P5psmGMt
ilpcnvAc1cTrq0NvmICX8SDxQdlg5E9Q/Ago93SoRBqentlGLGxSNdfO+h8y+JoD12079MQ3hRrw
b3EsPQlbOY0JoDgH0tbvND3g9vxel2pNIWPbAHPrim6uAPrSuEqtBRrvErKhWSSO+baKJCqcWevV
H36xqWLQQA+Sus3UCcKO0lbwm2+oMKvK3/oMgchAWnMyNZEitdIXJt/BVVgRkESXQoWLofhM4GFy
0Urs8MX2d/NhtD1iR6i58evs9+6nATk33HOALXN1jgntWhPyruI+GJqachjurCJws/LVnKl3StZL
LvAioQ1lNWWhIthNVCYW5deeuorOh9sImztwV06htdld0gd99sQnnKcS/u3EeTbKxZo+ISA3t0Mn
sAttVjb5Lx7pDrMDdlLDw8egghekCNuKFPBDOGgDm7XCHiucsS/qN+mn6exsIhFR3bzsDXisPg6X
2U+NBdQ5ybe214NHzRxr9ustDd2OvShQWBXqcKAOo29jS19tmjQAmlIoUxeo/FbDLLkfUTvVtBtf
7cto0OUKwidjfkjj+zZ9E25Ue983JhZ1DF3hOI/7LDHEcy26z0wKcqgGYM6Z4uVWdEJNgwIst1j1
bIodo5EDVamQ4x6UP9abHaPjOi5p1YIrBQJ0jG2oZWhdPpV01VNJ1j/OS3BrUcwPQqr2foP+ihWT
M2zQSWL7pxGR05ZOiI4kBsg575DhTy+Ud8YvEXli/xXe4Q7sEH8QMJOMXogRH8CB09B8IztwaTri
9FM3NkH2L+N+WthgqazQb+DSXJuBv7P913jxvVvYMtdLWcuScvJEfPB/od8/jDEBt8o/HVfr7wUJ
LtzWCp2gw1WG/2dfNANF9XvK5hzVzzk1v5v1YvsFl/YEdo9dgzT0QEqkOOw2XTxAGb/LZ46y+EWA
7J/dVTGfkh6qLELkjp4G/Sv8KqUdBhko0CGPnIVpWiLiyH5gumO5Qst2fLN6TCN0LZ+2D4Wj5kvg
mLJrHfvUPyOAVYoRAwX6xjsa6SZr0XbKDSS/M9EhuAeEvSowJZY2AdLBUxuHOPvP7z8YqTeMLDV1
eY6TDRxD1bS06Pp5tn5aChrYRPCKuMqatxETz9lJjqKNd8iaRcXVjxikGFvnoYDasB/2UFEH0t47
5n+86nFvJFwYd1gh/X41SvtM0jjSkooYikhkAjAAZyQ+143wC7Q0hg4HdzOPxTS4xUE3VbyTAYqA
vl+r3EawTKFjE9CHNjcD7Jsh2qu8D6YeV3FjphQRhSvbSF+gu6WymVJlbMSh7qQkYRd6OS8RqgSN
eKcvMw6kJ/o1x6aeDVjJEetWDRswiBXplQRAnj/87r9pAmML+ie9vW2d39tYOkhrw3VGHvpASbvT
xoeQtlwFS8ypodKbt8jUa9A3LGr/aBPZ1uYTBWTUw8c0cFmApz8tiDC70n95+c2u3l/ycsSFiRRz
wWjtl725i63JF/ze1X9WymEqmcJh4QH1QUghZFADRmTTaeiwsSRCOeYhS46KMj1LLyY7NWrc6Re1
ljbsOZCWIk89C9JPxAcfNz1Tsbzdl4gXi1/ZyShVP5gNk5UX745rH+4SWY03oWLm4VYd/Yngaioz
chJvQ71NBXnQ0aYIUaO0eUfRoPo5NXCuWRpnaAVyjPwKJdB3bEdhPFRtiHqyRs4nPA4LIJKmvWQH
1Dup/Kx+5EyOK6ByQK1Lb/+WVnHsrMR5tRWkV/rszdnjg3JNdz8lKoBM0jix+t8BgsUMYChEw9mX
1tcIWKNtoZbwO1ABvQ+VTCEP0WUAWbiQpSA6lIhUoWWumUz0yIeMDPCDQyu1gvnLhYvmCieqSfbA
IfZSnoTD0eZ3maVhgvwUYlgtOH79HPOBqXnfagX+V5K8kf+G+C1b7ewoMG7g+LzG2jkajJI1o8Dk
ka8oeQ4B/kM+xKr/6UA8AHYFM6d6Yd8q/XjBj+2Zts1hoIZ5b/fuhfpjwlihI8B/mvibmSRugC7r
jdIsqi1M3XOM5b2x/4eXC3nyDk1SvYR1i6IhR3kI+7Jmqht7otgJmyMYlaj7DV9XwN0vprhgsUsq
l6xT0sUQPBnV+qYPPKwGoG73fuwhDmwYubwzey1GhORQNZ6BuI1uNKO0oKkCnuy5RMbvUj9xO3R+
EO9PgeCraw01rjn+IKIdxwhswOUng3TwpULjMQkTw6Yr38+oL4U/PElv3RfMc5gI4vJReotjmOag
iGXh7C2efpA11Uqp2/SRf3q7/yGmcJX19FiT2MAPz35aiaI6Vrp2mKymmNJFrwMUojc7GUsoFL05
KnM0nD4TWt9urPOjugkNQZjq5OSxyFs28p47EP5xwnF+lfLdPd6Q78GgyboaEhaoD4PL63+qLihE
/3sRSBT+PARIkOqrvWxUO2YrsjyN1hfahtEor5nu6dI7ydKoMJza6Hd/491rFL5zzqeiVh6hD/iP
mz4VSTRRCjHCeZm1I7IA8RihHhQ4nD4IWYSU/4VZgh8sFySqfOxXka2XCTUv8DbTva/+3UaHp4qR
cM7cjIQPvbATjf+9geRS5eTJrrtOaFAPeu7trVzRcKhwFZ3kkaZCvV7vBq306fPnz0c0Jb8nn/+0
99JiNNC9jD5A11k/Z/qfRzzrNXZNB9KxcUQTMSQMZrpjZ0CHE/Hz7EPW1LnjMqHOkCTzdQ2PSpAo
BkHChQCmPxNHXGAs2SNC1PY+JQtDZCK5MpjoQt1wdqflf/LTlY94iWhms4DBpiIpe4VbVQ1XI3WG
JR+0HQElpRgrTjoVrRMLl1+jZpwo733tJR4lDlZBqVvxHXv7f9qX+NRTojfZNRKLeY/k8D2MWLkP
SAAAUGJ1hOSul53hWKoavzcMq91/m6n4DDTxcLT3Vfh1qXJ181oWtfoGn4r7vGu0Qj54oCbRZ3iC
gmtoSAcqz63UOAiR2xw6qZ7diHGEYgnMFQN0B2FzDSewjqS5MRYN9rtiHmowknEHYTojRWsIUhan
8t+Cm9rIzIpccmpMrU3TluJtvQiC5PIcG4NDEusk9h5yBxK4fWUaSfFQ3inu3yXq9ne7k4yjQ9Zl
Mbf7nkghzChr0LOZ7Ihvt+WFT8+Iv19EGDrzJphM4lKWBFA23po6Dq7vZZVS2vC8lFBqnjFP5esb
ZS5z5mykL3RaZ7onm4ApaL8sBV5ZDeexkBlgtSRmaXLr8fY5s7pbwFzZ2vGfAJuz7RIjlzZaYEj3
EOKfJ6Rp9gRI8dcPZ8i9nHHH1x9G+ODicTAF6kCto4GZ13natsoN1EtmCPDf8miL+HGX5k9Ec2Fi
x9/h5EGESxOougqGJrCc7FhPLcE3Ooa1Rpmf/o4K6p2QaUXPk0gM+ykGB2SxXw4HfYftUUKQXY1x
cEHl2LXODWZHB6ATbJ17P8R+eotemaYaDmlQrcKGn01IvKKUWvD9UzRMfVm0LQ3n7XakgpM5uNuO
RkkvLVAh/x2wx6lvXuRDg2mOpuRDPojbdjM8Z2G9h+KyVqoTjphKcUx64tMvsLv94pNO+LbmZHSt
AJitQi1lPCdLL0jEplW0YYHHrv9boH9QpqM+1ESTn7Ai0w/F5H0zTqwOYYH8AyMBV+jxblUFH1Rb
pIktqBFQXWwMQiTqaVsaOFCg7uBwivMTv0YARMHCTKrdRHOFSejMb8AMc/3zi3X9OyvzmSZlgR9f
dzfcnyWzqpEoVIAqKp8mHKjBOw5y7VKw2Ha+7hUhVhM6APRNLGO7SBUBxcvA3qgBggp/u8XLSd9g
b+2fLBmH0pvjhyepQ/rJo7y2lGS9BkDJpWEKVOggdANfmXcZslRlWS1ordnYm7g68ONzrRc0HGfH
fZzgmdW+2FIUgMlVQYTKDAnrgG7CJ/VmiPsM0JiB/7bmrfhBYFlQbDb8KP+LASOJOcvl6OBVawe9
t1sNwJiIOR6GUy5Tzw9uVOF7MzKILiAmYQjDClMrtBgCXu8PyBOO6hKmd9qminB63Bp9RTauX5PQ
bEiNFO7AtDs35CBw7PowiI3LDPBzoULNCOtmXKQL91bdL2dhNySp8tdYN5fQfpCNht2X6jACHyju
ZS248omVUtH4i44IcmEFb8LQ2/ghIjT9SSHl+IXZlUNN7DwWLgXTXag8sw1ImGqkHxMsGUouXkmX
dx61d8Au+GIg5hX1kLJ8FmeKQwT8r6Uc9i0NLF6Y312+RN71KOu7D+tdkLLRScCIpMbaflgX03vE
foZJK/OnBHQ1I3KOxQwJIZNJ86OXOmMii2sOd7l5+pctjURRnUIpkD+VV2z2EEZhtkZnimFfDwRd
5CgUUi6HTqI2oQkDu3+UwO5fP8Zx5IcxM2U78fp7Nb/092JlrzDXgVvc4ZwFAFoA0kLz5//2nxHx
5TEXNYuaHS+nl8ru6Z/A1GG8Uu2aqCERf8LLYJ4fmrwx0Z66u9e1hyxvNIluLGi31tdOy9IYq5zx
C/MBKTNarKhhVpxi2B6fTwc2J51VcELoQufnJZ2wlZF+IXK7ae2sW6WoLwDrfpM0LYQrAg19auq5
uca+UhM4FhDl6H6xWJY37WY635aMYgfgZgUOZHE1KUC97NPrvPonAYc7QxzCQIaTamRycTvhN6Vu
AeI1G9RhtWR1I/2hUx0Defog92K4LU3u9zuzz7AAAN+9TW5BJbYqh7cxS23qsfpFGE9DUF6IS+w2
N5SKJI82ohO1nDHtu0PpjoAe4IgIauJ5v9OLmNWABrcqIu1rL0JfW26YqYOko/5KWNVUuwIu6jOs
jQtrdkaIFMzLiMzvhbaR+NOlJCx+j0wt7CmDk8Cdf7uhH8DSU7L/yCBjs6K2U4NPyx9X5D3nc2BV
Mp9SgWj4/kqUJr90ylDF0wEAAzIgvrtECcQxjGv7uJtaNHHC1B0EDCOogKLlbbhRwfXbMya/3XlX
P4kkHGE8qnxCzholLvlgUkh1ufrU2fywXliQUAxrQbfR9jeLhZMJ8J82hpHvNhWPiFGBICEtySRK
mPCD4sQld1YvW9cj56MettiTNiF9a+RJjNnjS+ZdSFTdeC4kB4abrw02t87xkPfzD7Wb8PgETaBc
hWq9wKPONFY59Gf3G+VqI4lQGAVObNYniMH0RFq9ETsNB8vfr+jT5DZl5lFMr2C9zGOIWY02k8/H
Vv1m1NRGajSwYoTnJ5BEfgCd23LDOptia7onjdcuoyrgvxEpC5J+AxBaMFalfLC0TfdGsohBPHL1
YQpYEeM2rtma/JSdVDmQ19o5VavEoUw2tApXYnVvX9EUG6vXFLrS8kVtI/WYnt8SUZIyqqn57Iaj
Xs+rwP1MW6Rxx1rdC9te6gtrvaqsqtQDFW2QPkWUp6KhNpoE8b86PccGTFxCkYDW7Cbo/CP9xY8i
aDSILOH39TRJE7l0mDPEE9GjQhjU03mYKxYePdeKHIadY1of4nQSxHHPP6CbUf7Y3gdMi2Bmn8NE
vleV+nmc1RS/vfm9SbGWAQn8xTZFjyKNewtXbILVf6ro6I1rNV/jYkwRLztDEBykiCBdjAWf/RLs
oXGxHTipTGintKJ4hy76byFfVmuB+lv8ZZvm220oL7y/u7VUbByVJ2yCyu0ocrrsb61l/BWf85w6
0RiifSY2eOnCdmMJ/MlssIiUYWjURjFTzn95MaiuBN2sYxQacOgE5ox7Ymk5gPRNH3omjLnB31Ue
xUQ054ICB00rsH3lOqxZD1Uk50b669Nyqtgw/E8wbf2LUror4bDKKhgM9OQP/20GG4r4ngtMPuXC
kdzh/Y+XEA/0+hD2LlY6rLxtGVGhV34gKzdGbm+o399XcQW701sHd9jnHp2adTxizWsrE81bsgGq
KjY5rI2VuwdPswROrGy4LTNpLAWPDwOToJExkmW/MYzOafi7n1k8m2cax0dxD+JDGUFwPdMqCk3b
gj6+RYq3S1i+VIlaMzC8/RQu3Xfe6mbnHCA3EtthcGW49F0puzgd4CzhFtxMUzcDUDabT6M5NXTw
o4NBunFr2qnja6stoTMoUZl+4Tt5TjUR1xHhyXQPe4XabT0KIuvGQ/609jTB+MFru9PvpBgCLpUU
XjLqSireD78ZMKWg4Wrs+3RQUmgeV7hTXEyhRnkZwREwy07cQ/HNQi3eeMZazQiBcAsAA/Fj43I9
w0jvyfZSDj6gSVnYDA/3Yvln3Hk9cdBeK6fzna7hk6qy5BOtNOzNRfLV094ilmHfZNZyw/PVcksR
vZYlbfUMwKXJiymNxRcYYRpJw8Tc85NcIweRzdNLRe7jxfxlWKVh9YytDehZSZcRenUbZIsumOWz
W5ab2KKNwpOHcJZLMx9PoOdcOF49ybEgX1cfTZMy437lh2Fr59G4Y3Deqc/+N4hlX4qdGN3mWuNd
tpY2n/SLFKpa4JzFwnph69zUZKHPPJTvNhlrHLtpavaFF3A6FIui7bJdFUU7kEix+WNND8xNSXJO
QvobbdMyZrJ8Vk9Q72G5h+72xOpJ1ELOUkajnJE6oD0m3EIjA7JeCCbA50eAI4dVn2J/MoVRrQyh
J4lNb90LCKrraPB7xMJVZKNwHYEB9sTvI8SHsgD6EhbxGaZt2WZZcrtSL/UoTzR5DLbwcdZuqWdf
CsBo0Y6s0y/CW0e/yw/6HSZ3b8rkPHHNnc+g2eWHMxcWNE8KfJwUOx2ELSX11HZmm0AshadahbuI
3FEoAJLIMtaakh4PfxQe5/h3emWIn5lTFsCk3j1mHQARKK68r8BUmZHUt2/2RE0Gksy6lMgf2emA
sdJRINErw29UVYJ+0QThUE8HJxx8TO+ItIkNeGr9bJAASQgzm+Y5SO8onCV2FTGtRJQ8MeutqOYB
RFu/pGIXPjWtkT/yUR6Pu22383S0z6j3hxhAJn9gIYOBTjbxW3IZlZSII4FWUJiCQ70Y/y11yFxF
zc2kGMktTKIZtnhzia4xd9l6uLorFvEiO03dLcJ8P+/YV+UWeG1NhgXTkZ+1LmJmvCz0ciSRgn4o
Kk9o4QHGvgYYBYrqjN5Bt1AkfWslpSd583qG4TzUOlKBwsctVjhJXWkCuCfpm8ozWM7kSF37Lc7L
aXxhRlUlmNfzACzoOLsplOl0ByuFEkrsj5C0fjEq1keW2QeAqg/K+lcGZux07t9b8yKW8ev9FKnX
psi8TBRzK7yQ8s7tLdbZ9McPmX11W2nukhO7lXJFE/u6mCTAPnoBHKZMSG9G0ZNTRHoKAsqHQspL
KDKXVRePWf7fGrHYkRwiXfYa8GwxROjtIuIOrmZGJ2RD8gqdFVkHS/Y44Jfwm/e7TtLYfKifleHM
jtM4pmlGksiKLIIDw0GWmjdnWTZY3s79UPD2JkDz+r1E2/ij5/N1EUDaNfsFCwsm7wCrcWAZvzm9
q9m4BW9WFfyRTXXIcMK8pp1arQI1vwZ2pO5M2CDd9/wWOT6L2MEY1S/VH9ZiQe+gA7txLn5dAfb1
bSyvtd6oZAQeVs9jPIlABLKCKAri5hy51vrM3OhRKAHgVFVgRkUhykoLCGpRavJp8WCQvT+IzBFY
q2TR9UHd8PkBKkF9o5Nc1M5jnyk1Irj9KJ4IyquiqgS+W4VbKNFABVHg/dm8glD3cf1yxsW81P3g
THlB7X/GgVNLHo4c0SPXlznzFtVBnbkTEatbSLB4VDNfvhmbjGljuR1UsgHn/XHlawmCJtgTBVw1
WUTCvpfuqt6vBC2VTPDO8xIcpJJjanRNWxYGHEnFOHFrsu4L6s5he4FPEqIcyrxRl8mhTMzs+61F
AoGdCyGqNLMoVSCc2W5SBEYwqwrpkorOmigK1gIR2aoPBMbRwv2QRILe1pgdD1r+GVALIlBAP75C
VZzGYB2QjnLnMZRMhAxKWYsnLU6Mc5uskn8oe8xDYa6KFvP+u28UMLiCde1eL8HOOoBIBl5xkAGS
9Bz98WjXsBjL6eu9nag380fwbURdmEyql2rP51mjkcQ24Gqgbs0NwtQ35QZDW1wSjyfjjM02c/Ts
m/2spdKceEREhy4lriE8nWpYwi3s/keKA6wqJTwkkjq37QQLJhoITioorptt/IDrY4Z0C7/Qxxey
f+nsQ0TV7X3CCLiqpAaY/FX6hjvPzzctAapuXdoXPWqQZ9c2+k13YIb6BfcsSLTV4t1kw42V/XTN
RAMI0AB17mi+1q22JczSYEUviwD8GA+Mc8PiY6gQ02jTinTqxJjZEMCHLTWytAjGl4rQU8uv66PU
zHTwevW99LDYhTE/Oj78ILXwnB+23GGDDWspgb9GQnk8fjzczVyp8qJeq4cmD6D6ZqCZSo73G8Gu
5WW4ui7bAwFSAr1n7y7JjGcWY4HY+lOlH6u1vlly9vzHFjdYJdqgjAdsnUq1r/Tc7YxLUV1fi36/
vhsCYprPA3qhJDEotyRIKSSuYn0JQEDcx2BmazJQahGYwwy5U3JRC1kFUsPzehO1y9U3qXgyxT1o
jsxmr/hN6/RD9agPzShlrcYx1Doc1ijcN4mQY6DOu+NkQ1tXY2ZK/LpI6N5TZe/u4FMRScMNsdsJ
adKhTfo8hyxHotGT2wISHPVJ5CmsSDDfWS/GNg7Dstg9FypR4Le3bWCnTyQjRIrgol5nz2sLkV5u
Dq9y2F9F35G16mQoS1F2r3I0Je/BZjO/4LfqD3Ko8iB+r+KGoV9IBIIlmo/tSxiNJJ2Jzf8uws4d
4iZ2iH3Wuleidatfe2FvUVfBxQrb4n/hdYblpH693m4pNAKZncqzilu1AtrzX6oW8BXIeNnUu2SP
vAGFVvNYSHX1u0OaHakvVX6NqtiNrIlOq4b6ifeYgDFuxN7aTkSgMr5YD2UDCj86Kqg024P5Q2jV
zH9O7WMO38D3kypf+/IiDxlXMx+CI58enxtcLqVU+ZDNiyGb83cKhRYGQq2ZbTRmfu2HjzaMcOq/
lM9sAeHj8JQ5EF9j/1S5SBpGEL+sMT1GhLBkFpdLbF+oEKjyxvjXhBHiPSJybGOR1e4Ew41QZU2k
Mc+jRLecL4Au7SQdyigjICfQvOKrk4Yxwjui1k25rjHFBGx3H0kGA/gZ9mY01hUQugN5z71+PRN/
7H0+UwqnsHa0ujuaU//RvTieKO0F227EkUR+r8tvCBc4SRPLX0L4TYcf6g7yxKIboWJ+FxW6m3eH
WJ0o2p8yP38WgT1p3O5mzk5gTyQwXtLA0MMtkDapE/DYRbOc+H50SdCGpm2bFEwJkrcQKhKAv6VO
NFoQh41j9aafhvofEZVmtYHuCrDFvNkMA+Rc/wsV9DaZc5pCGNQcHDFBWeI3xKdirVoTvq1mCTJ/
fO8tWFX0H6062Q6nk04nrbA56H1CE3q5YydGZxoXpXIAIFkpKsP31ZsC1rg6qk2YygDAdhRd53PN
ksL84Zjz32pfcY4M3aYBVy2RA/vb2YW7Shzt1jx+hYaMZnqWXDRjyPAoEckAst0OSZq2iik6FeL9
/WGVFtfe7i3QV3QAGT1vKK7cAF4JEg33BcP1tj1N9SGp1CgcLTn+TV3zKhtGcNKfSAQ3nMvD/14u
hO47KzM7A+b6FvtlSkxgbCtEtS+3OK9yC24nO+Tl90kuzkgaUHNBQx7/SpbFnq/MLxP76n00iWso
7X4ZFoSzkz5xGK+/VgUf6hMvCFpEy21oO5Rrd+L83JNHB4vOi5+5BNWWV0ZiDtzqh484SjTMHoRu
m6SEECBjzw6uo9sRpIOP2+c5IVlhk3imd+qOF7Vp0idQAuStheckDIa8G4ojpiS6i1p9TEcpdsOf
pDihtGbSusUNlXeyD+hGx6yI7PNz9Fvg9t7V6xPKid6hjMI+Y6/ZsMSHptc9ftcBaD2J+lBQXgHQ
ahHSdTvI9ByYPrsOebkF9Zp+vQfwxNebxo5YqX7M1Iw1yujjns2Mk6PlmIb1eBHWr8KKAGEUXfAz
xweReO3XbpG1CYuVc34GxTyqyC+cdeDn0UwlBeDg8znDzLn/cLbFA/NSmE0V/UFYz8+Sd6wxgsgY
P5xvuv7f8f8nnspPt7iiPA2xm8jljnEbs/mUCPIuJgf5UJoeb+CcLyoOy6/p+zsAAA60ajNlHlVZ
hm6+nLAcZRUytMHZLoe9mt0lGGjs7FLHIMjlf9izDF2aLaXPjuoL9tR5SrWd2oglSpxAVsW4SprW
8y7VKdNSSiXNyjff4thDt3OO4CRm9n33yEtmVF4DI91rkrtO+K0HuCJ4+Fy3i0IASzcUCDAKJfG1
Tsd494kr8Engkn47nNKeR2APsUdK4GM2mTngi37mNOWalESotCgA1dSYsKaPIeHxeAMzoaPvoJe+
4FzJrGGnfnqSUUWE+hy92XBQ6xdnwCNet7GBF0WBsHbdLt86/BjOQD5CcIWO64xdWAP9DaM4NHmC
fNkmG0vaa5EGrCJuqEwgJalWgFOR5irJXd6aPoHgHRQpJ2pAImTGogXxe785d8oaJGXJwfeGgEEU
dr+3pk4cnQGAJ8EjFGXNo272Hy5b97ocD5qJrelgCxblIiuDXaiqobEOfAD89eluNNs6l10r5gk+
SO2HN28miUVnDmRYXMEbkxbVIBc3oqSiNbkWmwC01qY4XVaOcNTBjZ/LCoSewInXuSbt8ZowEvst
enfzMFIVqdmgjUOR7Us28EtY+HZaiNRY5/RFeE/oaoBdj/yN/cikEEKj9lnRJnUhmIAZyFWztrQ4
ZtmsNerzxGX/ICioYakZQithpQH7bDnqxBjsI+YVrP5b1rtuXdsQlZBSuS+zC4MQeL7h0rcSux74
0exGW7hlZFmS1buLGkl9sX6Zo3hpVv+91u3C0cdpraqTlcyTYuYBb7QRkTQomsE+aALfJBV9KKVy
EOSPGNezW0EaPksZg1ChEmc2F8YoKxI1KV64YwWQ3LaRS8SMAC4k3v+/E9oQFaQqvWZk7ddPk/m1
sFA3/HaYk1dm/4o3PKIh+auFnF+W03zfOJi+lqwDQS4n236XBETm3P9py1CAY/eU/ZIypxj8xGme
sBSx2b0YnVqPHSScVKRnolfAiekCHO1AvTcMPdBRwmA7gDCaS8qN7PqubmXoaQlCergRFQHS/Lti
g7grI+VlyfiGuzKMTsC5J1myqRkwYPENVaVL2VuDxdJEBokuFXwJIxlM9h+Ln6DkfcV6RW9+p8g9
dbGuPhw/Sl9XjPU++/Xd5ECBWKHm3SfNtYl3c/xwW2ru+V4/muh98J139aiv20D1bS8lt8njRWIp
Gv0bABN5bLPV8uv8pUHGVHEtIO0GXhHJr6eioV5FC30kEmDiHmWZwey01oYHTHWf+RfJW7ctKLI1
FJPFwj+wC4X15NQmANq4XyFkNT3kcCasY+0XzD6gJl6JM/0C6uSBD1UbDOAWJHDZGcXx09NqKYEj
Qe732qslubfvrB3UaNmvgOVnuAsYFs7HKnABeQ3cLC9Dre+klfSp59i2EjhdvqeU9i7mCRQ3M8w1
pKhV/VRQ7uR+wk6Jrz/jKcE8VpBn4Jj/ZKn7Zbf7EmuvRDsqf+aNuuqEQpgrGkilfNXM7VNhpnf6
9gSWRGVaQWehua0oU/hwPRlnNFcu/JIltgC9ddvUwwhecVjpFdH062sT5lbSqcBQdq0NBjS+tzPK
9HpdjTHRzGkyc1oPdhG/765pbKLgzgVtyLdM6B4YnLB6BqtZ0UdmGs8OepCWOEmEOrDetSl6ANyQ
Z+NsY5l/UG1qfIG1yh7xEP0ET0tCuXeXmmGEyH5xUlLr6yqOaIVSfdMejvEhdcAKqdIosTYmQ6iu
BT2UjJabbwCXa4Aiwn/4sTrydtj4uT9oz89CibeEDwP3D/IOJ806oafgmJiHd5PVYI7nlo1GLhdI
h3KtGBDc4R9xCij/KS95QegrY42g8n2FUT6YFgk/Rj55uBtwnes/ddCDM6+w7T47O3FpNtelh4hj
VT61Wvro2LEUq5KhtLDsbAZ9eLn3eQbU0SIZs2WZgajAUyX0CUwOw2dxWgtrLBOMoqTOc4mwKo0k
4AeYFffrqPomkM33BAcWjYXjRJm+Wp+XyCAQu4Z3VPAfXc/nRyNL5bklt7rkKFsm8yhjasAb95pk
riWqJ35/e8TaxJaFgRqSnvfh/WdvT3/qvojWZ1dHo5wFH9s2QGSC/tv0jwvrCEZe1QbwyB06KOiY
FO0bmlWJnf3Ecc8ewvqmocTN2bwaqQtYtwB5wQKBcZNKZKwqU2ii6TadLncz5w5dppNQ2tbzWO/t
SR+1YVtvjcMSvKkSPSaDJmfloPhpoGmd4ODvQJ1JLLN7pDwCRb0IRsb9cinaHIkEEmjUfZuab1Wh
QV95YGEZ5jagxOHqSrLy7h0XoleaCR+m0MtMcBg4q9oWgZ3m6/gOnFGTS4lAyUMvoQVofEHl9+Q9
zXEegrzPSP/ZZcc+h0zi7wusKnhuxZSXPtesLbwx9o1NZzv+65tOEZwys6ZHkeh98NepBhrHJf14
Gxq4l8ns5vzugSP61RsKBvOah+JvhsNJAhHLinLIfEgL0DYV9N8OOLlJVe3WdFQb5GaV+Y6a+cT3
igHr8aXp8zE5D8uyPXHgmc7l7Erbg5vzaTbBlpK0V3ePWjjgPusq3tgjX5Kdi+dtrCXX+io077hY
/xrwz3G/t4CaImpDyPj6lPncV+draLTxM6ksnmf2z+K7+VLkbTbu3RGCwCrQSeAfTfjv6fN/Gx8b
nxkgXVZhr6Q4Ko8LIJAeWnHDV4S6osdiEkGC0WjDiCu9xWEMPAgCLhoalsxNU1cSOxTkvbbvaczA
zX4WZVgetGsPh8g5mmTCgowLsOdQL4SBFQAABinGi9rtFrgm4z7TV0bpKYjp2EWAB22WegFRoSqQ
s/9/AYR61Km+OyN79rTuclLUuRwiarZfloI4gxfHvibk4VnTSYBah26zMpXtXP2E/cCsrYn0LZt7
OwXGYm1lweFzPekwyE3YUta9EwhNQkNcTNDWQomejeenwBqAUoo/kdIfBpRvcQpqn/3bRFD5TemD
RZlo82WTdRCU+eYRjLe+4LhhYWoq3s4TUC74Gq9TmOtDffEK9x43/SF0sPIEDtxpk/+GYSiDYwNp
HLfCiQcH4Ycv13MrVmLVaLBghujTk0EOm492MS5rjHwUY9tdOdzV+Wt2fSsEwmEyKCRzJX+BFjjt
Ws0sHaYozR5IZs7/s6edTIYzrlQQpeWImK7LEfqCUMLNjDDO7fx2JPVNU1/g7ctx3ZC87HefdAWF
CGbtkVn+6Gfy4zObWjOKUppJdCoh1vUVUkfKtyttBCoLO8Lasjj9Y+ymJGVgyDJIXSIjIDgiwl2f
yItId17vBXZN1E2i8lab1+8urRaQVawDCniIfX7aD301Yx/3s7/YLnuJziXK3YxkjO5Hae90vBUr
YMunmqr3/Tr/ebe4mhbCMaQ9jAB23NSmQhqe+bd7Y3mwymLjlszo8/xe8fYj35Ws0UfsqzfQrM2q
mDPfNO3h9WAGXo5SaD/HUIUFcx29zEnR0blDb2WSQcy1s1fZOjZyPIrS1VtBa6q7AhARqIAdSPkn
P0H45y4TVdTrXX7JFuS0zsQML+zAK2+Jl3rTXRi1Q/U1Z9VQfqEVBEwEJqd6oO1pyQJlj1CeqVX1
qlWY/y4EsxSmldlQhUPC2omTSjY3Gra0uy8UOmJ4EMttteUgcHEl637kw+D3FaAbkURoxj8ShSjU
WkeMDuYWllL9azUjF809EhSHkVHRqMh6qOGaldsZn7nCHoH44+G2ap3NB2Ro54oltaC/FMjPpR2H
n0K4zmtt7P5cSbR2g760DPljFQx/PXclZK1+yW8dhhaOONJ+DVx4JWC1Cd9n8InSUXTLPGAeNrjw
qFVrVg2KKTsag6lIvXBWVqgBOeA4H10j/wYpooNPZuUdVDUgcB4Rqcarr7x9balVVYr8SbivXCV+
ZX9FLJyEqhC58vJ0WK7+oXAHQY+qKAKbVNz8SQnMQQmSo1sg2xvCkkDI6F0yR6uwUWCgxbwzrpVd
6T6fT3RpVQcukLLCrbJu06U4OwOYa6QEXjvwZ4keP2f6qxyAS+S88lcrtVTOtWBNZPN0vyur1YcJ
y4mkswtx6+p7vwj3AaKS01qM+bLY0TrzRtCuu1swu/x6A7yg5WyKBpK/H/xzNNisaoBW3ka89G5O
VpFglBMHD7CnqJMObMIy1z+avc/XamxewQLCmsXJ00IU8VjykbXjp94zluAGL/Bbd//z0ZwryL9i
iwLBRIBfSEFNvzHS+DN23fL8fDZfsuYHgJ9ry8wVE9BlMO6pN5Q+nDHcOgXpphiDMVXXPJofiR57
jn5IjV+OytdufgP1qX/VUGWQs7EYA+C0G/BoN6tAtHmRFhphzcbOu6umzE+8QKN9sFp6Y/DCq2AH
Egw+LBvrSWULKHEOB32sy1IHMOouYMycKu5qmUyw40Hva9fNRzSVnBdsjPYn1tP/IKJ5CFlgTdlA
ojsmXPLIbOTD2T+il506nt/nD2wLDaS5JLuZQ82h7h4vTjx87KirDIQW3tcc0YUN/X23/7xYLlGI
Gm8PteO1mmSeTLhCfIHXc7wOXolYVU8sxJRk6lUy3xOhjNkbeDLdQltN0iGTpXLS1Vu0HXJ6nBu/
x0xRpLq2fM4i3czB6NyTuELB1w9n/sZQU2tOrryYwIcnYaWNGSHmDUrJ3Eqa2ThUgg42vy4k6fzk
wX3D2shTfkkHBzCEJji4+E10pEF9361CdlZQGHebRVA4aF5BpWkYA9wwcArw4MPerSGfk7FmmLzc
RS0vEHMtS7bCUneEHiF9p32CPxydlHNmN1eIvvuJQKP5SHzzb6veMIiaW3HPPmkTWtoq44rYKuMh
xp46xT46zPPeddnf4g/RrKb3aEFcI2pqj8+D0d0C0IdkqZ2WPPZ/G+KYMYmnYscBX3VD/jbn4Dc6
R4yLpI65bmtDwBs4bF+qfqyfh+5zP2YUTo/fDYPXHVTesgOY1CRHxnhAFFQ/qfQsXBUwq/MET06f
BoKBvSrNiUxt+w+6tNsvFrhX6Az+8vlZ33QgfyzLrumL3b6AK7hEtvDJpYdC6Ih7eHbVwx9lDxh3
pUAAOhvfX6kDnNQqNCkY2nGtMl/Wy5vGLPLq/5TCtrUDHTWKcNMYywkiIuHQMZggXvM11LVNh2iC
1JVDtm/mt8sYIX2j8NcE0QIYEbFn2GjCbkJ6RtqG9FqK3e7CigCXsucBhFcTcSMtqeT6Ohd+ApMQ
NN6G+EoAXErDXsU7JpnaSdM9eYnZs7lEQGm/VWIzmTKxRLOdIbzmsyZZlmUhWYfY+PqBMJnxBkew
cXpUDalpL0+uI8/ixENn3vls26shDi3DkFW9QKqSuij56QNHLeuRvQM3coxIjwPhVwSFcNU1rUkN
YnvpO3elzA+hkwwtKzgZt9oxVVxKx3cMyZZbDZkRywCOBkVQGiPK//HwL++NlphHVkh6HIv6DhtL
HbljCX4anJFysn97uuThP3aopvY2Z/rhaf7PQGUMeH28NQfE3xRKxG65XEBu4Qr8ENKzF5XLwz2G
J8oInX7mTZZJ9Lvf50615/Obu4rsK+uzYN9x3EFD6riKpWFZsxWZGc0JzB17Y34Brwm0nGr8eDbB
NyJgt7ceGlHSCehl6S0+27YLovkH9GKdrxss5MGmAI7mGeUQXUCqKGHYuCUpU4ULumcLikJX2zf+
M+gbP7tBOI+TVMlOy/fmJszK5pCMEI7RvudHE96/zSF4HwSOZL+gaeQunPdV88bGcbEUxJ0ef7gM
+aqMMJ2lehlsiwU7vrH7CURArmBWBk5ert9kMB3WoLB9nvbEbALJkiiI0JAPF8ZUUGBRrQblZoNZ
JrK8n40Ed6iz+SRw+VW8wSWYXSerwN9pVVmsEuEzybHEnWUmU3/RWE63ck+pPhvot21Qj8RKftS3
knA+XYNqBs/u7CaOJO+UCL6n1zjqcs6t3zjTzugS9c5sWZDuETqM1XM4H2E5ZQikim4tGrQa4MaN
zpnNRukqVqaTqZpc5FENZibU+Ib30jG7EQEw9PyRBObCNjejth04xeRHr4YYEGRZ6nC7gx4JwiKm
HxmJ/emQfCs17K1R4W6vdEN7YPZp5mbNvTPwi/4cWswTM1kZHQ9MGHLS9R2t5XIBUVHfZvxEmeJ/
uVz8RhPNQ5GcfMaUVo7BS3aixLl89MJCbnhvJCo42/9exoxo42qkP9Pw/jz9dsj8NCYg+QtrMapI
XoUYfQG2o/cKKyMpYFWwbAuGBZ1kccSwqmPFIMPSPevxNjpZzbGQgbTcN3SfOhtA90i63+coWye2
vWjMecmYk2ARHXx+LdjSWZ7BWQUB/T1ea/7gzbLMhG1Z5Su6XNpe8rtkhoosiGrbxTxwbp/FdwKY
pUuRaiGxRnOsBHQ13D1hL7RXVMtEhRX5FQmbY3QWTtsltxZ+WTgMEE67aptE9Gmzm4nwxJZw+jv+
lYfVBn7IX5bohLosCQjv7m0dNhHT4M1jND7VFX00ztYphLilA+5FyRqLHvYMK36lAi71/bJrAYqr
tiPhskCu+ifaMmXWQ0EcXXi/egHnCrhe9E7CpDeAdx+oQ8D9aF9X4xe2jmpowimUe43Sp5gur19v
aq5NbMH2HXanOrIyhKgiGSuGYCfWf5rsc5CXhKO8mVysGSJXgmxAb6SpDyfEbuwGraQdvelFehGS
mK2jsWIBxivmiRbesO9TBa5WSeoQrkzhMzZKWpop/AZv5qsnQ59QaHQkJzKChRD+orydH7y6nqZI
lPRD5O4URATpjcNDth+iZioyM+JPCHP76H2ikBpu26HZiLlL/vHQDpu4VVbB+/H3JPDpzcZyzhho
D2XqhUvsO7fIVdjua58jdq6b1At/udOl74sKoZ4v1dHh69oA8MbMdK5rV7xXiPBWmymaXj1yN4Yh
rN5jFuBRaFGCmmaGeL50We4rb0VgSsaEgSNPUhSuGYovrpQWZzAVkaXNlOqjiKgRkFWy3Mu5Vy0x
Z0dLf9HNco/SpoWikwerAnbrkFp9hm1s+3bCsNKdU4s3XazC2Vq2ER9yD/2OJPCmzo8Z74aKuUFp
iZEdiXVnpQ1L1E8mi35hTQK+ElLQNuNpxosyi+Jh9veYDN3LZHEv1/XrEtUwT2OUMQIQ42qSz3GK
9TwHeREqu5YsZHA4f2q7WHIQs+Z5x/eTdZwJUWKQVRa01uviuw/Ra/ZPKYYpmfIdRQfdW0PAa4LG
OJMYPfhhrN4VuUE/dWfI3kaaXdbt8SIXXqEXZfwWyjW2Nzlm9JB4T6qXidsW4PxwN8Vxys5x++bl
K+OgzAYKO2ZekrmTS2dUllPh7HCIvJCiqTTNr4oo48xgCHVPOggg/OVRTTFLWjFdvc7t1i6zpp/7
H5Cma1gn2BOh+8OFxqOhcp0jHTxXJBQZrF1Tz7dCxiOXtKE2KZllHQJ2AI3Q3/WIk+wPx4zl2y3G
OXfvAkCHV3a5VznPZpa408S94ZW7YNNhs+fiLIZQeivCSAqsb9yqb70hIZwGpntiLb7Q1dYdW57U
o3HJrL3cSqTX6m5KY7N5F/zR3Ep16GmDI+qiQJiv7IbP18tb141u7W/HZuUVcBvrEnDvfJI+VK7K
x0EQxrKk0LBRfk66Fwv2WZPPl9PcRLU7Xg5lH8ges61nlcmF3rtTnLhbenfxyu8B6ERClnfswK4/
FnJBV2pnr2iXArSeGSMqRZ22MgfhHqUFBoQ4fLO8s5J7Tkm+47vbeBW7K+H8mnG4nO8GVcUYfqZ+
elPFrBYa7H06GTPh0y5NcNUG5Pxe6UAGUkSpPeNmFitN2fgNdXK20s60Hc2mI+0VzF75WA2Vm4go
3HlufO+wxgmV1GEvwRvrJtF7RJ7WtBdYlS/OMBIxOsGTPNDhErGd81Cfu/eGDQexTq5MGmTz8Sxs
xVj6dUo3oQrvz8YaKKMMNUCnh99JMwFZgHab5fNQfcRSDFKu/f5cw+LHDbD8FtatFcH6ezsi+1vc
4OwbY3d+F9itk3wWqklXP32lS3gJvDfYhMjAQfIkX18xlQID4xF5bzwQIFghp8uaC64wZDPYjLWf
edXcGr+JAW4UhDjUBcxckkEfOyuqxG8x7hti7uiYYx71FkIC9KrzMzV96Ne96QCIwJvIp+zQTRiK
AycG4TmWP2VG4FTECXPCYv9PEC5oPXMsy4Gkaa61QAJilj89kQLIx8SjzSzVbI77w+11mEpwitz9
25Ek6tdilvVJTkjbyUFPKAi5anTmxTtCTKacDemJ9r9bceyXvbWcXmWPBOm/AsE1Io1fvdLwIBxa
ucynYf4absgxRyfczgzZB8fqP0Y//oaDNC9+SecawRoCgwcDHljDkHzay7GcJK1lSfu5QDh0Kxx+
whffmZiziCPEP9PD6zSdhAwpFMZlXVt66Sl/QMf8EhBnyqYtOsOEZhlatjAxl1H8h8Pcdv/00hSG
40kdK7XlNRkqaqe8oGz55fQK8Tjn2nmv4F25/c3/ApyezK/F7hj4wxz8jUjin/Cznv0vhWIhyZDC
74vk4fuGsxjt2vS8Tjgi8syI6XOXHtHUKbRba798wUAAxNnHwHyB2Zh+HOMywG3LDm/qDlm3RcPx
CzbpRhY22Pk+J27Ejx0Yx0blOQ4xL0mJ4d491/wj8/uZfgVzUJSXX+iHQu1y+iIs986YMAyAL8s4
T7p3HARS1WnYzX9nKAGxZon7UqI3eOajwJDlg9gXXTybPPaVX1XzwoaplOyh8O4wKHYGMF0tai24
3unrc3/Jm8oBcbIIsrqTYMr3hN0fia8scBDgm+FsJeW3fqOC6N+mlNThak34ARENFEMD9+3IH6X1
jLLO+4ojVPNO84YM5jP+Z+BPJnK4foa6BM7SzW8E52H3vdZADxcdDyFi439IjwXSZ+1uCaMhcnRW
Fdq6KECyU3izI9rwDhhTzhfJGDS39w0cfkmI7Ekr06ZfwvSmWDPDDvPk41xBYcJf25spSbeK3AFc
oGEv2QHAIClILg+O8nFkCLuYlnirjtfP59ARc8h9s8qvY5yaifkce6PK2/UQHnYZTjuz1+mKaG2f
WybAtHbg3lfhsos4g3kWYhCluJ3dEdj95cpjt86Ue/VY914FoxyjIDJRKT8HwPlW1PG2cnEP5pZh
h3rtORUkMOUzhP4Hj1T3jEkRzgiX/asXb1x5EBm+QYaIBsM8ELeGmYfxrkERlk9FEPPQ78ct0Pg+
Ynt7Sj25XFCQjA2LN8CHwEcEv0fiqoHs1PNqMK/nuqEhdjRVbe++RihRImFGbTn4pppR6jtRmlAd
1+ZVskaqw3enNCaObfATK7T8zWqJu5SCg+SdiEcdZPS0R+W18Nyeye+GA+xsaSKRHkcIbrUEZgMH
Lk1d4TDzpcrG3VQETI5T63xve+ahJO+uSLUpPyWbBTahc7H/Gdw7Q69dvTXjMmbUms1gy8umN+JO
ZrS0MEDVCwPOWKLg19uoEthVjG94Ojcm17qtcMeTse+7hl/ewTZ0Qw1vkL7NiimlS7BYRDSYr+Oy
bdyJmLTQ0M7mbYFFh4Z2JhvaTTl9m53fyyO8wyjhRpsxRy6ZoxVGyZ7CQFWMXOSoe64yEVuiqkWu
MJcsNEZGCz7JrN4Mr63Y6zXv3STB2yy20xTayiXkQZxowOigZZz53Au4q7Zx62lnKBUmA9dQfTS2
4QCy6+tqGszq8q+Idugq342mMXiWVrBcGDoZKtxxXtHB9KQJ8jL/HG4kx4sr8kIgscjLQ+5zEKFW
1YZ+8/2alsDOep41ogHKZnZ/nrZyiMEwbMyRYOVLRVBLCIMa8Q+IRNmJh5UpCnaMH6RutnKj1tTC
T7w+KLPGOpnYmABQ6JXeJZEVyoreUOftxQicHSmlLGwCMcWHVlOiO7v+HHc6P0TplKzV6RdawmC2
T1JgrfvFpgfI1cAZxmKF15iVAdgj7oVo0qWQ2hEwP6JsCrHvL6Qni4cElEPzIzraB8MJyQODwvmY
SOP6ziyjy8JdPMh+zsMPOvk4ZRHWo7LoT2d9PhLR0+rvwrD6aS0G71HSxO9l58CZ9Z2VE/Wt8zsQ
xbkvAd656XSWpnPM1aOgnQ+VBXzB0sRaBREoOxhJ+kfn0MBKLjGRkIieXwlVNEUiKIYsrrbGKEmH
V3MaHzebQGC3w7KBziBmCh6HiOoj/t6+U6xJ2AlqF87C/wxHwNlMCf6KKgrk+Uuc0SrWIl09UsUt
np87dX5WtfQBMmurwuaCWUDNCu2iLgGwLderXK2ZNaYWelnUhLpLCJULBfW8P4GqjsQL2DG3cq4i
k3es1mm07nyHMcupqEkuktIV0GHWjVkdwMyoFdM+aTXqpJYTBFLeBQ+ZGLTUwtakEAGcTaakNzrH
V1Vfg+W+VztPwsTBwdYc7ykAI60TWj0z4kj/7dqHAYd8ijSmlXtGg6BnqfbEGw0c5pLk4hm2iN9k
3iXf6nQTeWHjSMKVWDiNN5nkuw6xvNoZqCOav2O+0BPuTcduh5+A78FJ+hmtWr6IMjBGPKbq7Kwl
lwXpYi6/BWEYN26lKjGCLCDZB4AFgNg8jVN6kT3mnoxTRe61A2ypQWnbpsxz1TCVllgD2utVDzxx
XJvttpqgNt4BDbpruhU4SeLIW8Bt5ip9pA7eaIO/+tmmfBA30Dp81OQifYfcKJzl/TEQij6b7bMA
dqlIb0fj/gbNgmdcbKNls783JdpTZ1SC8XiTks+hKpoZmWMj7FEPJo4WDrp3Eo/gfYpB3tem9O8r
QKaSelm+ChaMpYjqzWrMtVfqZyxAa5IYh2JhmFKXicED6zJQQ5wyyeH8oduKJoMpMFoPCwOq4PND
VJc3NWLH+Puh3Iwa9/KiaCTLXBHY76QpHHo/oz9bnFZbeedB1nGx1cNF0hUeOUMr2Vi29b4EfJcc
J4Vo+aLLzkP6bdS9uWg42awxVZCMQC360dZ93V2tKjO36MRsjXpVexffauCA1zQjqsqOsvXsYKkx
ZVBiYku+xcFKH4n9bPyj4Dy3V28tS7nv48m9lsFAXPVS+vEjUO121uarpGlFdWIbhSS6DI2cqYr2
06Da0glq0Ot76sSMopDNFqmzB+uqwuo9vcLpp1EpAJtxyCve493Fq4o2tDtUFfQm+9jPVpRUOYOz
pHMIYbFRkddpFGC62kODKnvhOxBaWFquLVS14HaMycWqB9T9htzDHnPUVQxdfJH3sz0yOwAuOpVc
tjsI43KVQV7pApqiYTEbYG/ctDmnKyoex4HXEGC0UqUrNOwG0sMLs1TAOLMiLhyW8KrfGpZmRgab
hPcaYv7fyY6crgMk4jXTE5oIrsEbGn1xhCKcYSCk6iSvbado9oERQs4IO66uLcBIsl9stGbRlrdJ
shOilGrB+ZJ74EkHNaz18ahsj5lPJfg31J/POURSRo2dRQoBIw/ZgiEtaVCeFJkgceZ4jRNsIIXT
pk39dzRgKRBeXNpSpoCVhqjvIFX/SMyQjdE1jhFNRn7TaSkJUtL7RzSVqvZeY5cDT7udUqL3VpaL
0jN/EVU+4hLBlpS7jKvOnglRb2HAobM0c8xEQkoE2zqUmL9eGYu2HTJ2fmFimyuvRSLg0Ob7Y+uz
fLBQKd0YGunuqD90UaN4cgVe1n94e/qCpQ1JzUFZE6AqH8kLw50MxIlIZbmpjj1r8ciEzF/+AMIz
CNWrnxjfjnw9mzejDOLDZZLVqIub49nrb9ZCwZ4ckLCvH/jzgTCZjWX0T1Dz4mmwVn6FpXEPf0lj
EWZtYTsIV0AMYD6sfKtCGhJdxZVXbviJc9nQC/DYS0XGTasxWbU4gq+sJAwGxK2vJeVjz1289w+M
hoe1ndPYakTH5tVRXBiMOWT+wOOrZGJo0/o4rHzSlFjhrlmc39HprJU3H2VQ3i14Mx+zPQO7Sguf
rzCnGieNXw41nXhvj/D9AdoYwtfj785IVLxbyWb1cVhEGkvYcBJ28iJ1e0fONKcYiWrfM8eFlFhC
YOJFQ75HYOooBzzT/rtol7pVPVOpkX9IwH8TY/YTWQzjVMHuSfbCPz3Vy0IfvV6qBYlF/vjRp+S+
Ob3mAB8MIEztjWCZyMvi7K3ylS02sGy3U6MtiVeibNomkUcHl0czoxn0KmGjXfvo2uPmZIDoj/A6
7NWr1ddp59Nx8xdAYxp9+3FrCoWxk90WK40uKe10ImPPjtNbXXWXJytN7vmmi5d9yXaV6k3oztyD
kLmfWK+Ej4UunDVSGsAY+Rb/JUS0sKCtj45Q2JzlShP0iEqnASAU02s1uJ3NlRHvK90YUkq/tdv2
MI4R5P2JI4WZXz9PQ6AOBy3nzcHh6UF+FRarH6eUR326kB43WciRDFhFV4qh0Y0FZose73Gqy3Lz
rsjipvA9pR0RrBrkByhNkgGjEoiFoQwvfeiYsz3NhPOciMgvMfSD6BCezqTHtGIiRiJhcv0wxVrS
hb1oI+9FNTcruuSmjyUJco2e7116gBsdEoTSTQzfvZzhzKgL2rEnX1YTpzRrTGbp1gQLk5it+uKU
eoMykD9mM3xnG6aE+3zkgueoIkTxa5uB9QLCrvCyxLuPUymHr9AVztZYHPxO/KHzlPg4qJMZGiy/
0XTZa5Nhr1+G4fTaYlAzXgfqF1LNvvBevzatep1ND0Mu5w3uXFDQqSVRTE8hgYyDfpAqQiRc2iup
L7ZbLeaPJmSEoYOuheqdWdsYBQK62Pr/E0r7j9DJmkERbtpXUrI0z2XaNy2cfLVEQ2Nx50D7WG7g
UwT4dbGr1GkDtmn1a5FXPmfZ6kLjK8MKMMlcbnTC7xNqlCJVGRl1HbLD8vT7/1AcfDMtr6js2z0x
2sfuyOge2mpZ1ZgCAhQY5B9u4exnyk03xaY/hlVslFGJAMzv3ACD70/HRYN0Bk5esyqp8E3wptC7
qrk1NlqAllUgIQasYinOMbP4mGZkIwgC6jWNx8nRndp7VXsY5XQuj6e/Fqd2I2ESAL/+7MdFRggX
vCFpgH/HmhSvufGRO724NU+oCPGEAXJIGZLZTqRAR0OMSGJJo3L2wHyQs3UuXxQmiQdtrejderQ6
NCVnD7+bwGVQx/uIis4w4wTIp362PKnUnx2t2n/mtBd3Khnu4SHiWDLUIrMrBcMT3PTtItzYFHPJ
Ce0gtQG5cTsCshOfipR7zTC9TD2cJel24FncrY4cfQqy3ALxBL/T2v4BcNUiUmfdmyHmFiIarVll
hkHTl3M72U9JoM7P4ql5otVttK5eazb1+lsY9853fKHz7JSDJ5vWM7IcVOubFQdBKT9hrne9atll
FwdlX6z7nOtr5+S11g8bXNYjpH1zBpAaKE45On2fN16/WLIJGrZ/xmQBSqe/Z+HGuewdFG8h4pa/
tqzfB9YNsvDwjgQycoVX3+atvhWlBB8rgyR1GHtaIv1EXNw/eFLvPIgu47mXFGWpZcz11gHPL56r
v1dNjB8Kkn6Ftc2kXH2MMhnEYso49H887LtHalezC1ePEFNbwb72V4QtzORwDg8aySFgGr2wn5ia
e0Pvp4IqKrvsgWkoCWWH+amwPAtQKG/CAvaxysKmv8NkZholk5bbQd1+OFEoEPFYt1Ipcg88wgLq
M9/ZMluC3VGoNc5tgLk76l1HL4D507NkAWRIKXy51wSRApDLgvK0/yLSRRmbAO978HMk3Vm/Tfiz
kSC7oFq//iIPFUOV+GDfcJYSkVClLt5vbYoCgQXMY+F/fwU6s1oT/Ju2XqwdnYYmAN4BhQ81odX5
f+PFrxIx3ha0KcSjmJfyRK/JrenS5MLTq631RuzuW7SFlMEatNu5B/R6x/i+51Wf58ygBkGyhFch
3j4jFKSVnr9/ihBykSIMRKuk4pg1bnvtSKRQ4SMzY6ysNpGN2E3tKOkmxVpIkrc3MNb/RPYkKyx7
Ruur8CAeRchYkSMFT/xFM/QOiAucgYmFs7NHdWOoZtcIvWcw4KUuPj3azzBH7HGzjhqGupXFaWrQ
0yc5IsNpCSypuO4Y7pAnDgXdDnYlS0mCQoTJbbGxRRCojbMlYjH8Ge7BYyn9mtFiSYZGejmVyIMB
X2UfXUFkB3w4ctfZWGeHSNFxkenbIERniiyQ7nUaNVR8wMzgd0UzntnixCtOcDedIRqBNFibrxB2
EPqlUsZjXFnnH/kksxvvN1QlBGgjR0Nmi2CfFOX1bamVIVzqF0AunRyLG8eWt3k2DcMDsN3Yi4pO
WA4L1y0ZGwxOnTnFujD5sv5qcJyzWkrma9gn5NtqY6mSfODtdDAZwmQXeyGSGzclg0YNqO27cciz
pfd/d62xLWGYcDQwn6zyZa8MJNaVvQKfiA1ekGeOAXn+8sFgL14f5z45y2oaXLlCoFFNn69BqCgD
aHNnh3JAY5WVwxxPDN6RRS4C3Dxc+AJZ/MXI+Y5MCmspDp1fiH8pgel1hUIyDUoPJPapc0rrIEkY
hfqkMm9w+hJk336Iq/5xPh+ZLnOw9d9p9XSgAOHjcf+QctucLiIQCILQ+WBzL58ABOusT2ftB0v+
f4E3bNbN8NmQCXrZBIx5W8lSbIOujmLU0PuqAbtUwrCZIGm7NxPQepUEbVpgl/0jo7p6x8Es0+MH
yP5fMGNVGVlifmp5fxWRhkvWuIh6KNIqooToBYfaxZRarAQ3+rBhgP3dzdarxYF+wK35nWPB3HBI
akZU1sSwkBsJKZa5qzGI6xOnbrnbhK0Znfa1ozAAfhKQlhWS8N+woq6UlCTQ/W+BM7lN+VFFzR/a
P2yeP6m5YhEs+wy5WK7M7twpJIxIiCcpheH5wWmKX8VbONS4eCqXwxkIedI+zqDgEMaPF8in8Ijb
96arOnDFpg7DKx3CNCRhXvo0QQRFiqc4Fz7+b81lbVj6jpPy1rQKcT5ELJ0cAoCXSaMIouE1G+Cs
5b9p5CWQueMEAWhlu9hrk4X+ACKSld7+ZpZY0cBfynFOkPwWYZpXuoLh5czX0WeFoKL90PToCqDf
5vzQ4c7aicPA89mqc17E/7crxAA1lwnO+6qYFx7AN1Le9CXN86mw0L7hPTmNMfhKh1z/nPCyuoAT
6k1fsiXT95A+RITyd5g4M8raIWyvl3ZsHCELXlkEnXgVeIYffsIB3QuGnrthMbLwAEBuiJthZBce
rkDt4KISdlXgs0l9vla6nnHmqHeTtSG8bx1AYD61AGjrZKNwrZDOMu8/2NSSSczPoBApVvFWKH2b
mgOrwmoXDPnB1W3lH+t+SWcWl+AI7WWfYdgRjz4NKj75ym2RdaX+zYA1Qb9PmWW49rh+1GilhSn2
e8k276uoSSf0lrB8w3GZKM5d2bbsB3+3rqunosp4aXVWkkYZEEnsQMIw4vNRQFNFsbcFjbGD1aog
XgHm/EDv6UIwsLmF0q6yy7hOyg2eoM9NnWRdmUiz6cMm9aK3dyT67A+Z9bi8DXHD/NkfxN+u/TuC
Nk20GLPnqhTXB8jwngc3u45ElEm01YH0IFzaaE3JZ/BcyKK779fio+XItAlv1yBwaAEI5pcEMypm
6YbHbSOAuo+fvmGhQk1lS9GuKXDsZDSXBAvCkQX3VnptaIbXR1J34fImGi6b8pUcL6PUFwF4RvMj
3YeHruBwBoFDebZAXiemUX6anQTucsxejAwU5Z949AGWCbhuK7okuMVEJ0XlS8Gm26e2FyqETkmF
hEyUhUfeHhUoQ0B4nmBmjXnluazlnRPjKJ+FVgmdmU2oDuONv6eyHu0PeO1LWedrVynswLsTjZD2
l1JsYhNo+7q8SANMtH6PBZ0bEbLPW3IfWQVdoUbU3gl9cyRJoETPmxpHpKR7fxZPX4aJe3M9F6QQ
X/g3c6bg/07HHfLB78gJb8AQq+bUADSXN1jx34QY+2gzEh5RN3KhurCcGFIafp4oeUo2UE/LWMzg
BdGJP76gWQrl/2cTNSDxUb7Aw5WubAfZt9R6wwOU+tUFK5oPd4od90/wJk+V8bO7sVmf8GNg0IcV
3eDsadB6oKdiPi+/jdtKWKcuG8KMmmLYHISa0UizYXm9EgTVMTX8qEefkr/C0lSe+O2Md4bh7zdG
u5ninwdKMHiLsHJUOYdu4ORP4AwKO1/3BbHL4LvFXdM7nPs67Gnsy0iJfr90lacQZ3MSP2e894ko
lCC1VbR4Tnpd5RGgV/WVzLR8EedyOKJYZsXUDIbDmpAslGJyxDoIocJXgAFFd1k9EPLIdPhqqj6G
S3JBi+J0EZdPoWEkkYLc33o0YSXQFAUZPGUXdjpmvVeufW86/SEXMo6Ul6ne9cIyDla1Ud/SbuwR
Jl7u5vwnX55oUnTPlP84rKyo+hMNiENlogJDojl4stoEw52iu7La0gXWHNUN3dIKvoMSuRa/HMcK
biLI8i0KZMN3lqvbPR9e+oHsx9/2aK9jlCrvDCjfr+ObwPg8shAesDCVjmhV4PR4VktxKVeidNOz
YgkGQiNqSkPJb/jzZjmTAsNlf1Obqu1igCK5xOmmKV6RyNRGY3y1IF3Tn0IPDjSd0xPA+1fdnD7x
jSSWAMtEkBAza06E/o3R5BlOc51dP0YWlA4z6FXVgt1perM/HlkrTjdUgYZ7gN0rbqqd6yi096qS
A84pKm1ThEbK9eC8nvFIkY1rHzkPYu4WpD4CP/tmgqg0JMoYU3ZsTNzTpz1UXyYAmh0nwWap1VxW
LrhdUYNIvi0G/n2P9fIQqjYnwCJxm60zI/CJMd2ql67l0MZAoZSABE2uRW6W59zMCUn+0MtlPcXS
X6Tdk5wamKLnSGEMZNfPtuBBrX0S229Zjviy1mQ1XArhAGg2NQmd+QIV02pjnpFHiOz1xmmMa+Rx
F+4PsYo6EcThuXV6qy2o4QKkZucOVMXKV0QSHoHjd6pGlnKDbZ2QCE1C8W5aZNKWwl6SZgNt1nMN
zjVZozDRF4r4Wq9CqQsx+DA6nyobwkhQ9plmR/OIGHCXV/+G5HmieQtfI33jf/U7u9sqxyt8HMTo
KjIOPafokZFv71TdX4E0IE3pJQRoLSN2OI3vU5CavFZcVzE3OnB8CU3DkdS1YSQRPlfPXe304WE0
zjcRMdy7UMUrbrxVgmoAS3iZPfcqrMWW/PWkYaj2sBE1zVHM87wiwToJX8blxQltKof4UofUUHIe
XMwrWsGI/vmHs2JFrWoposk++bKrNSvV1w6HWuPNu+f0nplnS0Xl5DqZN8LagQRKSloeG3FppR1d
hHJZy2TR1Itohjw9ngXhm8Myrf7tH4XyMH82yAlUG5/SwrETCIW1D8PuJL4/2aPKWhzuZduNOKKu
wrc00wxhpGZEBRFr9k9cyK41i09N4t5Z7oh4i5gP/sKfgp5QzOD75qvvbUmiridzfVa7Qm5ZDclH
YKb7gJNJ6dtz/7TjjeqHMTNUoBI+AJ4mFixl5KQtm0gtR8pCUBjHZN2292bRhG6XFBry7ajYIO9L
Qcr40gSS/T4VmdWnrSMEwCAOUpGH5QWpsATvtrzlpLR9JLdKU/mZSExpkhJCYbNs2gr86sgNfRfG
bXSL6uForRB21QOa1NfEsxb6jg3WwglW4Mc6oIyPVliTYeMoRFVQSYwbNWAHVKCYDhofhvDzumyB
3KIcACJ9F2MlHJ2/cYpaskp08YrQ+T196QWN8onBwpUobtOBZ4qXRH/YLrzyqJqsYA7YcWx5cmBW
60qDFxdb2H1T9rCdZ29It71t15sdZktiaS33ZNe4W3qofFyCkq24WpkOtIqHXOlgC3rOvLZJHJbN
lfVk+kj7HM6i5o0QkACQGVWIQORuq8IsQizRTQlJ+x/ieQZZkUZj11fGlF39PI66+KdRAzRN0GVU
gQk2JvFvU625ly2EzYzpJDDNjTwuXKvcoyRxpHKNgFmAIjgyq7wj2zE40kIdR4q/GDzpJn+76q2v
voUPKZaWjKPHbcxl69kvc/7EHiCScT2B2C/FI0aLun+6devsX2TI0U5QrMEB7GEhCCwMIAUz7PKe
l22eoTS21ohQfov0/x1xXQXHtV9PB7N4YNaeMh8aAlEIc/Sk56gLZbW5NolvYZiSoZYAneTsHoRG
3MDR46kEmNJ/wpAc1NDQmRSoMxaADghFxjeHHVJLBRWJWu7VgDHZpwaHQHk4aeSdKcn4yb1CP2iK
KTDP32WZAzM8p47VmyEcvpCJpJK/AckGxgaa6gpy08htSIWJY0Kilse01YpwMd4k5nlddhL6wbor
QH6hAZoMF9fKkm1xuK8Z/peZ3yuxI8at0N+h9yqorEzO6Dvk0dQR/PrFeEWdt3oJyxjHcSR6rPLq
R+jLA8jh/KTyddjOyJpBX1RBgsdsGC/zw1hGChucLiGnwqrIs9OAsPpKN1w8uPR48fbosGMiLLPJ
cU1OjfYJKJgseo0Pmlesje06C/K+xGKhEiWsTSrewdCoQVSs/ggjHyodKp9hAFAMVYcyanoAcR+G
hz1cnF27T3OsVJ6l4u9tAyfjd0z10ZF09fi0C4HhxtrQwpVeO6VwS/rtKD2/kn0ZcDxpTpi7jqwl
anHCIohFrQ4tNY5p5L5UoWXA72wf3eAX5hTBifz3eWESBEVifDW7m5dhu1WLmIVttX9mG7DsPTne
BBAEhiS3lFyi9N+KNCZINpSAG5uH5ERuTBFjCXaV6+pycxpdHu/hvmPfZKuMMDNC+P+ZzR/4Gt7u
TncBAvAwJYuQB5t6zWnnYlTSe7IrCjDedNPY5SbTAiCIHuMRngb6ACSXypQn75WyEftM8Jk/IIiE
tq3ifSbzakAXbXqjNDHWq7b5MQGboSkdDh2oJW59DHMZQ6QiG/o+sHxWg2rl5OGf+jTK7CE3tAxN
tZ/vOeX6zFZQxUhSYp3hjUhbtIm1kW/oWwYMbp9ABhGiuL7M7Lskhzrg28D3rWf62WxAT2A8zfJi
izCZ+ERVUytKhKNfQB32cKOfM808UQYam+k0Ax2/dizN35F9/71d/6eF1sq7efl2BHAUOiuu3Qij
hM4WIw6Z7zp3/jLaOffuwzLgun8cHOUyP3PSifG7FviMHymAUEL621jrJCmf8/U6vR+fV6UA+SOL
7Z5jfJgrDXTXsue18dG56b2EPT7IDZetT/MOefYfb9xx/GSpBl5oso/ksJfDRv71VM2wdX6SUQS4
va67NvRXsSUrxv2XiNrVpc2o2HW8LmmT4l9Tc7oaiiLo+SgUOTgofPLOGTyV6R3SDokxLgdEXQOW
ZCvWxlePi/C4tEknEK0xyQ5BWbyQy94b6oBpjoIZx6l2Ris637tODRZzsDdOihqXy5ljJW2Vq5yU
PriwKL6cv0xrbq62C4eswZo0/ZaRsnxggoke2K7nNpGPF5Y0dmh2sT06bFMHDXkmoQt9Ajfvh2G1
3nfazF5KwhK/AVs+7q3KGhMVdL2zUnTUlKD4yMp1B1pBizbtPvlxFPImkfFnq/xpZzhwVmhM7J7u
DAF6+aKMI7sV+qhHb/kbojkfeYG9s3P6iD1TuNobZbE21dIGY6aYinbAIT0MlIPjBvC6bn9PPfLC
O0hDibUhn9NZvs6z7Y3OZkc0Jr50kOjF4Wa4e9/M16pUtifJ6M3hYKns1PQfMjZEpceQC8dZ/7/F
kKzx8x6supFlavv0Ep2nr8pvUWO/iatNu3fDFGmPBjql/lXvtRBtRu+RmVHApQJ5x1wsPGTdEC/4
Q2SA8y2WjxKWwQIaJvDsXohDTg4TDxQ6lkT9fmyvjyMckkXmfOnBNmxD/soPW6DG65Z3x+1y/kOm
gn/dCsHx5HVLzs9XL2iL6oZ1LYyl2mUM2rq+pNtOcdyjLsJxkJlLC71QqNad6GZXQ9xbcFuPlMet
mWhyBYBl4y7r0KkAN6HmXoUC5mY3HNp2BGGNzpVw8nfRMhLHIXcFsY6ZggwXwDh5nSfCdrIu9cqp
v3YqgG9Fn7Vka41dw8M4Q2EjtuUinGAoBZA3dK0vjw23b/SLaNfbc8OWqGS4/pfnqvhvzXk0+vZ+
L34SWi6kWIViSedMGqc8ssgA2lQFrArRT02Sm20eptVGGm7sKaVn2BfEskP0F25+J23zYff8EMcw
ZfOtqZO5xN6jey+6+uJXUK1c2DlnDWnfufNf5MMisSbGou/gaJQZLHng4TrlaW4m7xA+5A9lJVaY
BL+5Wwr0sbrzmYLWJxI6Cjc5iNMVoVN9zTYJOqG9d8lgG28vc51lYlDojA5PqLlzxEOFDCL7ZdgZ
JVi1qIui/wWpQkHCdkc0a12bkZuYpCtWzoCo/7SqepamfTmfSU6kdNv1lgwqb2orOi2lxGojCkAM
Cau5YKwxcOlIfQCCXA0IEhGJESNtj/v0CzG3hsGzbcj+E7VCGiPDUxS1/x4umzam5XrU1T6I4awT
1z3jOAkHmDRbPhr8OKUPUPam7+KwlPGFBexdzESoFSFvW/glj0iEuCqTIoihxGl+sIpjejdOiv73
tJS6a8YX+9hPYCFAH1cKlP67NazPBkPR0gtlwJhJ8E4zwzucdEpLtxw3boOgUwwhgjRslg16BtRW
Ie24KOH7PKA0Ps6wGAvZUXrhA33tOntFeX0qZSrgC0QA5spPhSIUk20COS3vh1gn2X7yDZDoiqWy
AOoVluh17AOSITDR8elSl6RW4nYYGi1ceae5k4icIHnRA6TMLK1eEwv5c+hMjdSgyrw9qF+V7l3W
lYyBFQJZOTLeGOlYiBlAC8RRhzrZ7PT9YiS2b9CDNpsG0NcynxFROdK8dddEZpxJ/5EeV+Ya6E+Y
OGcnry+RLUEallDPs7fYphcia1/zNzAdO3DnV1t2k+7dDWxOSvSTpi1ccLTn2oXPOjLGabPAxJqW
/nQrBUIVWCb7eVvPU8SgHAamOBmLOMoFid2Vf/Oj4CRc5cBn9b8p+taQLbVN988Wt4YrJtvyTpQf
ORykyNCZYNkwwgLTpy5e122w0PS/x5b7fx6sWUDS6MHUhWTs11NVLP0r//ZAjpaGSYnkYGSxEoRA
M+BZ7SCoWfRMRpG/puAEwX+BTA6LXTe+JO8qJyi0Fa12GCMzJxxMVphW9+DBohXFoukvuG5Vr+/j
EQz1mOyuM3mCEipjQ4y/w++o4Mul4zxyNZkMBD5rUa2xCFB5Z6DcUHHxJvsFH2yS8A7Lr0dAoJRy
G6KllQlVXPosjMd1Nx4VYeV01l2M4m4G4xlWbPlL4jVVHz8Gd+S5esKzmCQWPdcte8n8L2ICZCvp
f0CxRymDyxdrWXLb/QYJLUEtw/5lsr+AMshfFsezQIIAWaqPKqIhiY+ighpIKE5zPSM7bN0/WtYz
hK6Q59a2rvb+AeAQ45bNtTtfEtUeRITV5r3NmDbHd3tS516sjBco2s9dTmaQtwJI80T1ZLcIMO1h
ql4GLkI1CsF8gbOnB34k+lLg3XGc19IjsK2UE9CW5n3NI002/HOO8nRgw3sVTBlpwbQgjQ4rl62c
8YiDg+V4+wipWkfJUqIhstAk3GvB3VCwdaXQvXDmCp31albxNZLeho1nVaPkeXKJhW1idpaiPwff
yRa8/tmgpBYTSugD28k7agqDG73KqIzBiSMVvjplgwNIYyx6y1wUfiEb6GSF3Rp97KEfUWGj+ADR
9oVvXmSGnofWBtjJH0XzWAwPUAnasIfVA6d2/ew4poxnlqJtfPQPTyreA1WHtq5uROx9M9PmjH85
Bn11voYLJQrN8Pi6ZbcWkk8DJQ+0ZqUpgThTSMfCQDcbgb4XQuYAzsQ57CirkHJctKSFY+/22TT0
NhE7nHSmhJlSyBzUw1e16RcpR4fOYWK570R5vqJb19vweK1LXMVaecgkktqBpAj3b40Fyr9Id/AH
KRJ3jYAFQiowdz4ZAVQIomgqr1PQFJNxNO7FOF74XIaO3sm1MSDunTQU/fBoF95+W3LmgLBpPl7O
cAeT03ilOsNhHQsqG7gbFPK0Zh+Q+7jWvJbKBSkrTJCkdrCOSLsVVMrdCpa7f7q1ttlNUz/QBUTo
aZKx08P5uLsExFP62W7ln3uq2ALPkIKhyG6dYqhm+FBuWTIm/zXXWYFNaoagqSIyINL3uPU33Iq6
gSZCMANKaqlkbaqy7l9OGNnzEQtF3dndE3sfK6cQdgMkHlLH8qdV6ags3kYfrfT/6rf7LdgOHnfd
qHrOZkvbeF0btlOt+zXsRAaxaFCywD75rdQhQzV4XbnebRD0UgaTPrVbcrtuhVqpwCU1lIXdPLmF
oeamtEKHwRMb9h/yBE2zeMOy4voG9qUUaK0xNb447senPLk/zgqHS33s+fLv8cprd6APD8A0VZVg
7L0JN0qLwLZflVxAgHQFr/O46bhhnIuHb4sgCaLnPiyRjjjWaTZhDpz4BpJ8SUYgw5Hzdl3rlNYv
JhVdrZI9/CMaw7CFqY6mX0uHKST1hGLXfpSMaqpMSbDudiNxFU8fZSe7Ca74mDFFqQRtgM8EMz7f
z22qLhz/DWBMDL5W98JWUTlim1wxFIL5Cn+QlTOK1PpHVgwqrcNlHZglyCE9iFhilpE6s9irG/9J
OLgboaymXkpgK99kRwAJN/v0hP8dVu6naxvVx54np6d99XwmP1ShyEtEVK9Z1EZHgAQYpT2Sw3Ek
ksQmsBZKs45IAI+I2ClNpgnNwgz4Rx+4lQDKeoq22HOoy1AHkPCbS63LZAWxUW72crWl8FvtCJYl
q4oq+gBWxklQLE76yYGmq8pKs3OQxvlhUkeQcn2YL4qI5F6nTZkZHPyOza6NhGvuB9gY3sFlC5ka
arBO11oS0TvcSvvs6E/+8fp+col7gskeDjABY9p3JYdZKVXPDFJBkVTyHTI8zuQmLvvXojOpKSAs
yX0wKYq/4TEcAT8oNwFQFLPYd3GMcos8CCVTJFbDBB0Yn1lulBftKHarADFF6xmv5LpOh8UzWHN/
vLp6bl7r3MDrfutKpZpkUVCVc+nt8qV59Yf/WU+HkTz1sTrFvDNErvWhbqjAASOVbg+wA70TKXeh
uxLNF3S1wg3ICcJxYXNcA6tZzFmGo1kkOu+zO/vo+nTbKrAFnR/t7vMXC1imEMDPc0BP7orElUxW
jnWYhQ9+jvUby9RGN0F+5AeUccTigAh4oMEuB8hTuOJ1LDCzZoA04/ndzvodUX7PqzI11h+Ir+pG
VgtOVS7pEgqu1cVdgxjMqzzgGdyG4Xlhm4fwnUIOugoQ+ifPaA6GkWnG/tTrRvWO7CXfqxALa81a
Ox93LvUaVBQfklkHOidKlCiDARoTZ7sQnyIb5n0CTpF2w2Dqv2rf+FksDjnj4qWvi0dEaHyKBCcK
Z77VOcEPTGIBm/YxYRiVNO1O460mGOt6FV20DUS+JBq2ViUrBIbPURwq/7jkneTkPp8gDBP8CvMS
iTnsGRegZusq5dJMUzIXYhdHxdSi1BXYpIqPJvJH893JjSQtJOEwu1WEWtJFrtgnyDJvdDI0Cbc2
X51hoERe6cYPUtfVdWCFW/lEv0oq5IHd+ZvBbxPzLuRft6wmSUe4nOmrzsTJ/6arVXBpBjXwy891
1vctFRVk7AJK7+lEkOEBFsB4N9lhIukXTzuP4nIhN+tsXxrNKKh9fUCNeBhLzPTiSRQIp3TwoZOz
wijCJwMY/gRT4tJFrhPuJ6IC6NPIM4rJ6IQbqVnMcvW58A+ePdvl+vxW2cTMERHF1fGWCIdl46yV
vKhr6ZWV+6mMC9MB0Qz9MOVpd9DKhH9Mt3xTc85DbZ2ctJq4h9dgzJEuZOzdAAOVm8fxc+kI2fW7
t+fVDxIi4PzQ56yi+87C7kJ7F8YzhvNe2R9Qax2FDuuutIbnoGP+p4cfYn4CsmtNiefFtGFyKQ2o
68eAQT7NGir8sy2Ejduhawxc56kgt+4NiiLKmbkOAapUjrBzilKfAjW5wE2Tw8zUw5gcGii9SYMm
ZUA3IAsTr3dv441gsQ8g+8rVykc2OydxxJ4E45dnc9s+3oU/+bSYYUS3qv7cpbNIsg6rMTkhbvgP
QHqw3SRr+RH37lw2yLNEyQ+QgfGfNEdtX32AnHLp4AXSmyN1Q44jKce7pjiNWgx0WBSdaIntsrrk
Ys2+8wQ1VUh+mgioqg0BRQKIDNQKW8c9nUnSP1LX0J4vHCeY7PCzREq4krEtXrXwT+NfuFD5SngN
xP/nt6EIDHykzzP/qIWY2o1bwi/l7NI2i7ghbj7/iLPPXcxodMU1EoR4mhbvZ9UgSDuRQqiPEaHG
NA82uSnZ4bPl3ROHE9Hoa1o/SupVCmwTeJqivzBI4dCQ5xozGy+40tb7V56pGfCDxUQn2qrdXEOn
5zZ3NX/VP8H6O6Fyk/X+YDv7eQYa8/7rBNHYuvwg+qS1+PtidCYHDiKJKz2HlmB/wBNnApVWLwxQ
y5FpatHSbv5GUqwYX7qcKFqyNd0kdoDjFfVKt0cjqVBRHAdihCClkqPg+Q6G/J35C5mo9v2hH1Gz
txhyJLYd37FwA24RdINRwrM3wgiC34iU/6lPKBw+sp+xCBbI4/XzbjnZ4qB6jnfLSy0e9eoXi/vS
f9gSsaJmYYM9RdO5Jdv+qERBMxbEQlvMDGHfbYVk2qS8Jy0TfLNF00UbSeIjvk+b1VXc2wNgFKsk
r5KBesIrmjU3Sk73dDNZq7aUfHyO14WttJu9erksUTw8uVzm7ACi77g35VQBt0EjlPVTK6biW5MI
sdWus4eSfq1zp8OF8C59NL6x13jvgbGRWRBxrAiZxM5j7hD8dk8nDHmmjVrZ7q40KL1UmkNIp9tB
NCqax2hDdWgRgQOTmuW6kQnmLKCb4y+kGtL3e+p08DnCK3QpPYBFGfePlRrxmGXHBCrnbHAxwRx+
aStRUrwAMh2YfUsLA7NGVLzELcyFUaKqUq0N/19GFt1/CLz1QHcOrTs6mCrJ//RXjUg4vsc0U2h7
MK5VwpPtGC396bvPCHGWd4rdc43apEZkGxdGdp+ZOsnnx4Oy/Dekk+dGFrXcu94fTppksd7RMwAC
kwLBSyxiitdC0pZKGHTJaFR0NYeDpVV6/i2n0iQMd34E1mOXHco0+nTx5CCmsgSzCamX5q3cdDZi
L8J+RxodjgfeuuzVa8aFhf/XsPebGOGo9MeMweuoqsoh6VrTDWvN/nUjOvNa7VFhAD9L4y4nDJTn
HqDHlhC/A8UI0Na6Y0DhiNEXyu7ezIFs7v4WpIPbDhTeFF8gS6SI2GrOYGyIp77sBFaHoaIfq49S
Lnf2ODSvL4i7NsHUp3qerxu3MD/Xab34P5Ukx2YdS+cz41SpZPVhsmXjKiMq4fiVTXXTBz2+wf8u
U10JOBaty27i+OIh4tG54OTOFPmdvQsA+q/t1MYJcRYZk3QErDloRmq921dqgZeO5IEvQlV2m7ta
aLYml6gE1CuN+qxUdqSXKPWG7Av8qaZooyZ5hkxVKnE2TqZsTgnlElL68Mm6CdZR6zsRiWWRw2Aq
+mzHylY7HvlCi0gPmkFv1G5MjCp4MVVrox3hmd5tB3jY+cJqRwheoPJ8/20Z441H6WRm8g12zM84
Q7yVXfUjAB/4wSrbGBz22t9pd39X22neTw3TQ2eaiampn+oz8J4+OY6YwQZ5bbQJ7c1d+uROC5rr
bmSZljQ3YDQSOyVxu7nWzd5RM/s9W5gCiWWZfoQm7nqcnfjhOH5lj/I8I3aizfHXQB2GU/jPJFHr
LbsO/mT6EMcN+d0lKHLo1YrkX5DRt3WPawPa1iu/yAZXwUwlefoSKqTI2PfY1q0Ywde/4NQi3wMB
ozw94hBkGXousvhEfVuCTEi2faW1IHMchZFKNNzw06fknITY+TRX+deykVWe74GlUMFE/VzbxroK
TCTKYU5mHuq0OUFvpDinRZJQMqlIy1aU++7qyV5NrjnwplLFh8FsgBNsPaZz1EXr2+BqdsI+SNEM
yKfAngYVu6YeViRKiTZmfVN9gcnt2zINolBjfAWgubIkKYSueFRq70L+g+RuFLs4vsGkZW2RDu99
SXpMMy6HfjYpPu+KKasQYfq3HnskOA/guC/1ovuYfYy3M8VVt+FCs34SZpuGntwFwzmnZaiBgvtk
GSBo6wZFoMTEO0AZmF8piW8p9h77HVhfZ7XtyjlwU0ghKKA9px5iHT8+VoDWGceojcOGTfJ52Xsu
9KQcSGJ5d3MPsb4xc05qY9EBxsICGYh4dd+nx0Y6zNh/SYJqL7XVl2ek64XdGe7wLnrk5eGVYZ3o
oypaQ4ylBMW6d5fseW6jNEDHQa6455bThiaE+K3sJZmtCGJGreyID0N7yyEKzCTukcJ33WL3a6fB
ogD61sF8TQx1/44Aba4937PVwxXzqvhLzm7e6SdLFGOTCoqBLpQynE8WL+zLDa3ekja5IwxUC4xX
YEoiASUCUyhvhZ/Qgvlo9DcjCVAot3CHX4a7y41z9ypWsySukQM4LVBJXpN+YMw2tE++mNWSulKE
dn11Y58L8N34A+3Ic3vxTGq7y74PGx9fdkVpBdm3fE4+vTEDNsmOBJQgM6ro9T5rK9PzgAAGIKNN
CtjFaOKV5wlk59lLkAIDNQf/uW86/OH30WmPopUk4xs3gNc6a0jNaVaA1FaPCgCIrmLMIf7hXFfp
/PdFlXcDtov9VoB2RLYL4vCAEjjGge0C1Wht3o59rQaazxZnaJ/y5lHCL/EQdt65RjelKWrozB40
8ydy1XcuIELyvT+oqjA5NI70GtVnNZv+01CejrZt+vnny3qQzb4/9nxku4cEtn+DtSXZsQSSVO4r
/eYxfDxxXI3Dudo2ZylBxRgKJFfjnsGu9Wugf18LSDrzMHHc2Bdsen5D8UCi3ame7RD2Xx6xOHDc
+yQuzTBn1lYqvWlWVRulAqRLnfK4i8TQAvD51OgqF2m3Y2VNGCWo6SD7y0SLPmXx6qc9Os1696Fj
grlPCuAAj2GxsEmK2Bym4lwxp5MwcfCup00rNPpz46NHPh8a475o4+rseVl39R9JnZTk4Mqu27PQ
HnwgLrmLQIeHDejXQ4FzDsxraZzGio+ayH9RWi1dII7bzSXdLEsHKd9d8213qaj3fSHkveR5deMV
k2I6ZnG08oDmskkx70NCtbVFsyy1r0/dQNTgWUj7ojoEKtjRjhixUSfgP1Yu4MIyBEn4Wf147XqG
EHgx9VC3S9UEa/BBZuoeJERlhivMVW4PJpFlAE1dV5wKAxvubsla8B0MBN4uRPYVEEG0SeJS5MOD
NcHMEHibuRIHaTsvv5U1Ak7rnEa55fOjbs45A5QQaxzAy/BGe542LkDLx1kADKrJGoR62jklsu9f
3IWTon2tY9htIdIdb/Bxf+ntzqJRQN6jBxfE84Lj8/v5w8MHN5tra8EO8FpSiEhigdWybrQdV80V
T8jA+kIjVjBRdBPTbJsmE/UJVDRlYEcrsRmk/6bbTeQb69oqhv3lVYW8dwsrgIyL6PqCkONAYSO9
pYoaVu1KqJHPJHedNsUkBY0Gb8MM9GcayuD3I7927XmATe4MvF/f59sVXcC0dHotc7TsRAelyeni
obCXtwo3fpzM6fVMHqp35lA9O9kTuWA2F4JOrP16dhuJQ6imOlfZ+2DPSSh0KCMVST0YX8S/cYcK
bKvf4RFiaKBEf9zYR3rrtF34PNnTpPvCeRYjEUkhklhJ9nQ/x93T315lNQA5S/rMqWRJqUZRZj7c
JqGol541DQGuI+UK9Cs0E/cFlWZyWW81ydkWoPTHibrv5JkP6+t8nYQCW+mvXGigQ4c8PfByuAmS
/Cjjak5KQdxVcoLg5zvyrT5nagRZiQDyEAJVEWwtrPo/QCEpRkmOMDm0Tnj47jrmveAnqw7BnpXY
3yjRIHzmIXSx7YlB+B3iMVruRYF3SXYTjrz1dBK6lGp99NLx6Cj1Frn5s5Lzzg210RXP9DqudNBN
kCr0c8l7UeqUcmDWbPL1UdVwyOVnodWhu/tqzE+GVdamJD1qC0wVG26l4mBmv7VqJZw7rK3jVGsk
CpcEdrc8t3gOyw43THqeYyiYMhU/cTkFgiRqaINpfjIyg3MUQ+XQJK5js01KrvCc5Mgw7R9Ywn7Z
U4b9uGfDvk5m+xX7oiBoUntOYM7KkJQxm+zUBIyi11o/5aSsshfft+NcZLD+oo1wVG8/02LrfOso
3ReUV1lHjfuc52C884xeNYHwutCE4o1uxKlABrrvjNLh1MM9gMjRBlZoqGyiWPCM6LtlSS3PLayA
3zNqSsyeJ+djkGFqzWZRs6kgH34vpD83xIR7BtX08wrET9Q3Cv15AYNfhYxN62KGwoh6VRZ0V3BC
qAUoSGPKcvrzxRVA6xIFYZTAPE/GCb8ojm8h6vLX1t7CMtmIztQkTgeyoEH1ZosNxulqTB8EkXfL
Iezp+aSbfvvkNU1dSDNXJ4szCNnmO54wu7h0zTf5yE3XgJROX48uwtnWeNuVYkhoHkNHATNwRX2i
KWVmTL1gmk/iUVphlmnq8UTfWEauGt8WT1qiwa+U8vm6pjlVVUwTb5E6Ki/FG1KxcZ6orajZvwWZ
DBm9rmurY0hBxzybwWai+lXH6BaIbkOYVaVOshJbviudbqr21d3ytkFB3g0y6u/fy6RgcP2bNY36
iee1FMLofRX7uIQfuHXaONih1SR3kXeyB/uLHbYeKVcASqcimR7PF9fwUaW7+6B1gNQG5ghWZaKK
ml8adRO7mKC0T5LxplEUEXLle2kyl3GVsO3Gtqevt7/+mJtKGF5GQigXysqi0LAEBLqbQrTzmpRZ
9GCr6A2ZheO1drxICuNG/XmmrlfbJ0EMXXheB7jdQ3kgdbkYVC+WpLvmDv2cib19jdCzZYh5gpjN
3MvD2yHKme6KzRm4Fwon/VoHiHrvUgfSvzXurRyjV+Ea74E9SJ5AQSoZgz+VqENwHGHIxB8B7soP
48rdcGcXhPTBJS4pYERBO8t2dbtLiF2Mnljc1ybLD8+i/zSb3YKapR1GmfKDF6pjeELDydcsO18c
yV6sov0EZqRCJqw/DMpNARjPVEksFKCaE4q6y9xUSSEDElV8uXmlRB1m7tcVUOCPFUm2LOLHSbd5
xclWDtYg9xZ6P/3hU2ueJIJluw5uQhd57xeknXzgH0Ez0ZYOk086neBiKWZbNfEZbFtYF/1T3oQ8
LZXWk7bWoVGljYbvEGS+ri4vr14BgmoUpQNUoqsj4egIzUOBEQq0agrgEkd6WI1bG7V4hXvmsvgx
bAiZuEXa/xHM6Jga3bGRl67LW5NasQ6pGGRbrcduUQvWm3/wY4ACEshPF6XyArlLHdYqv0650vLi
j52QpWbDaE44zDiH/WWeX8sPUiOeGNN0dLecDsOIkaetj5PUdIq+lGYPZrJFmHpXozAM4IYoNWS3
RuPoz9b6Ka3kWZMrvUHKSlnUUmlKq+5omglsDdp3PQ+r0b8uDNLDbiwqwxYOCfx7B/hOTLeL0QzC
4cpruMLTO6AKcL6OEXPUfIr6B2EIQfuFSUDjkQ5OvWbUxdPVsCscjPPfvKhltBQtNe/6WGKixpgt
VfLIRHW2aefuoVwvm9NKCpOjPlRj8lDprVNZcGEpfGnKjjVyd2+kiF2HB+7Eo0x2sOqpoRjPu/9D
sSsX7CsV0Nvsxz1G+/ubiPn/q7SnHoc7+xF+hUiJwVcmbgf3ZGhh3OtdoDlN+QDGkHcK/5l0MjUq
z/GGT03Wr3fPfTxYqfXBH4Xn52uiBk0Ch8be90wZcxqJnkFXrFb8orDgCTdyXMzvG3jvunYfy/El
Hp4cM+dtbOY8wyfNYFZndmlgn/GM+OJgQeBXGPFq9CCNAOaUBczJe0TUI5siXD0bvDYEvpi3JRZM
ljkxa8NWCtZh0fzuzKISDClzvHxA6RmTLPDuoZBEdnopcACgfiU/bh1yUiEQ9bSNxOXngiMrtpLU
kiqWnv+S7WWYDwyC6MqN0d0sKSRQa6kbHM7sIGNqsLx92W6JhZzSCRcpBwF1UsVL/n2cjkCZi0k2
glroC435wtjH6izSYh5hgvrTns3Y2+Fmk1StWpVj/2X9QMTNSndK05xt/kPPc1YErs8hr0uag4FH
xT30z95ohpDboJGzJ/ICBx59C2SFRQUmSsj/Nuy0PRGpEPjrd7JNu3HfHE5di2wOLM2i4eXeFGaL
YOi3wJdO9j+bvkcpjKKLmz59uBhyWBC6ppiOnaIPf3T0wL5By+oV+4SnWf/ypgB4SNCIV/P4vnG8
Ua7E/c8ipVZOklvPZaWSad6MUaLVE4DrsalQgIRsHpWlu0StO7bSe1tY+NUx5KBdFLuNdgdPXJAT
xexY1hhzU3FIj5fMrcEx685/N8acELh4vH8e53n4gLG6zo7NYuu0/ZAZV3l26g+BBG1AA+GEUQ6R
lBxU+HLv+W42638MKsqRTNbHSuExsFm8g+3UzwF3zBj41oWRpGxeeA1YmLNHF68PvtIgkW+XGVRv
3TDvwVoy8+GtUkO4ppqQN5UMZc4u5RoeCL1+IOx4v1ZSfiH0NLB/pRdVoQOyf08NR3tChNHwOtbR
yrP3MRtRXgFh0kbiJIZerJVzZch08IZDotWFBuYydNotQjnEkgTOWxjzyId3IsQ7tIr/5pGemXEg
je1wr7Tgjp9CmEQxikBXbR4jbSp/EFJugx47lO4fHuWr3iaAuhodR4v+gR204KVNbV/vIM3tVj+f
lAaovUfaMlT1PaapwAsG5CH4E43NSJXSiVYhmtD5/FKq9bLbdDXISqa4TNTFai7antKW/2BwsS4M
c/jvFVfshAxVpk1ug5SsLDX6ikBTiKp7kC8pWtVVB++di46KaS5SMBKTGbQ5t4UqnJ5EIAgXojNs
TCkVQYs8val8LU3MYn8SverRRex/q2hwWZ+G+sUTlAGBfFlfF0tnvDnv4uLdqAkm2L2+UMX0t9BP
k9FkoLcURz0Nu0w83ZtnjmOvn6cvthtl27oiGP9g/oavVS38I9jPsyHul6pHSG8WkPBIox318Nz8
rjutTc+XWYwD21EXMp2p+cAL+ZEKKKMriAIYvsgo/6tetdOcQEHwYKS9ZV0FGxPPMemLtp/cBYuZ
L59cEtMfC6tT804e2ZvJU1aLl9J/fpWe8COBDK3k9DsZ3Deaz+dG3li3gwlqaZX0QG2u1LYhdTf7
bidk2DYwRmF9BSHxrSJAS5a0YHcM+qqKVwH5ilQ4CQKGEw5DlxsB5wXZ9rz5cNS6Qe4QGskysggr
vLbHTJaFP6Kbws0wNBp57Cdk2l7AVaaDhhO79bbO0+6jvaokVfNy+iO7FBul0mlPF+0Um9vGOK1E
JmfYPb9NIm2GfWJIlfVYc2CGKoEIfAe/xzAAAlGTzqEZPsO3mdSpZ/OU1bKVviCGB0NtPmLhNpXI
lLdFzeDK7DSULyrEQN9f5J348mV1tONUyxTtzsqZNfylCXFjOMrXOBl92xk0FHWuC7BaVGoX0xy9
dxl6KSNDiV0+KPUXmFYAFD2SOipX/OqHCtMuwV3hCPnscjSyuRlU0LtL7AP5Qt1wKzxP1H+hSDCi
zeeS+9Yzk5+/MVNmIcO0vlffI5nETHaQkh4sAh0Djv+0HERRGt2MZPjQsZFN5Umb52rpO9v4wFjK
GZmwdx6mEzM+gU64hxTqgHat52qaGdNi9iE1HJCeY4NAdB0foFmsyD7vcn60xDZL/vACeCdU5P3D
yu6H0+SoeFHYDjjJHvhAoAu2mMxMYggLC7rn8J0ZRqGH2fqdTg3xGbWYG353E4W3ePPizDymJUH2
nEmInZpU8tf6htpq4BmR/Sw+1k/Ew6YITKYoj2sOsJ8qa+9FjcXjBvbQiSay1YsI5v3ti7eM16ut
s2Zaz83EINo4WUZnARliv5OpwGtTaB+qJCp+cpIUl1jWSFnWhpvIRU/1CMYgFQrSDg4Vm0mNoPbJ
nOwI5kfJ5Aex6kqa8qPKSvpo4xM8Ix6wI7i6rW/n7J6rm2FilgJsnY76zUklgrCr9knzzZfdLARW
sJsHBb4Z9pY7d5XL6FQ0kTdW3LtlEvxl4/OPseKtZ8sNVWowFUfDhg1Ge7qswm3JztGR3hsozLPc
kHbjNHIog6A3xW5LwcfCnjGd/7DSHLxLj6FfvTQNYDXMcTUfZlXnjvUIPJIKYoMHi4WyW0QYwSFB
bz/UywecrIaPSYtAR++K1l2Ag0TpF7PN8D98RYv4X0OXMzVhUu2dhiInn8pFbE1hhVoR9hfSmjGP
M6GPH7ZxFIrVSpR5HeL2l5bUKE+XkMaHmm2IxEOupyw2diUBtYIIBQHq4RlVGH8IIHCzYfFBJIIo
McdMsu6Rm8hq81VKLHQLKiJBxbxhUMDIIi3V8KcZz1HcX6ve7GbJQtJQcSyX+q8m1s1Z1Phb3AA9
/GIEAuzHOJkU0bwZUID8QRjsDzQDmxI3BJ17lfglaMQJe/f9dxTQm5BCD2O5w2bL8j+twAOx5yOe
x/xDNaCPw+gDVKC09ji3aJWrTGUS+4LSbWCYgLV+AD/Kz4hvCYgIlhQyp3CO5Z1RumdsNynoeyrk
K3+uIapnfEL/GPgHUyNS1UjPBLiah7yJMRw1JkLgDDxOpoCpO52+ClKmqSdjHmfkVKBNDrTuny8i
rJhISJPvCTVHCfEsI+tUV50IsHU3k0koV2gB0oPwqug0DYaY8f8gmOa+OmJQhcXlyI61sW53ZPff
MlQYJ2HY/rhWkjB683QK8Ek01XKDBpPTCdNdrfqxJqKUn7dUUDzLv6TA0XRJOC06leRMPvfmaWzu
SYgGHtvvzzMCzxMJoXxHf7+VoQCjX0ZFO2yjunR1F14N4yIvS3bcH4maDYYPzzedXyZNRU2GT/gw
j8ylS5aYX5UvAJn7RVclSh7grtNEC3aFj8RAqRkrTtNtz7iyBWcWA40dyPyB4EysDZ9dtenZ1Iwv
DvnAOicZvV4uw8sTowjj6jGR2vnGnavry2s5e1E8xjlkQ0bWxrxjqmW3gDxHBtgZFt0WqiqWYcsC
mgKs3XQyGZGkizmDeV6ciV2/9fZTfVjoMcgCHSpSW+9QnX1mToaBoOXT1avQPExtJS/MKAAFiBrb
4P6CrIoAxcbCaT2NR3Pd7KjUlq2D9clD4JY9YW2mtvo/SRsVwqx/5GJJpLaaMu3UBV98aRuJI8z1
+O8j6lGXlNyLCMymJggPDNtS1DtI4jKFhc6H9UyVaBuClwLss8b2t5NWA52nTMAdp3KVqnj1rvwY
kfIEEWYmJUQWa4cpTJN1grqtLuHzsLYCZWAH8vLn2WcEncoofmCQ7ht20b4hf2nk35uOYWkk7v7p
91F59NdUpGeVirqnqvEBUeOMrCrqCFB37FHHLDWKQTpNuon/5Sfz1Vn+k9rwwh07XffR1/5JK68A
fV6RHAlSD65vum2kAAi/BQKSWLvoCXuhzQ/Emx9NMjP8jCh6eoJfdzg35CsuPHxgGXGjS4TeaabN
umwctmitDxkQL5Y2u+0ZTgNe+jN5HVOvVMRmlSe1p/mLQ2a8JsGojnXDxkcibtUtiIurvwEsNfQ3
1rZh450Je5PR/EXhQh4YCpqgfShX7EWZ799DWpOE2Gd0smDg3gIWgM+pRF4Qj4uaPKBbsNMeSMZX
K3+AsJPf12wRKbsKQM+9S8UcdMZ2QKoyMw1sR7fMlE7NOSeVs2Y+Ms6S5VUKHUkHcGVUDyWlODOA
WOV1jEzm77nbrer8yx+Nqd3yzglugARrMoLDcn/K2RxUfWikLyb1tPyggQ9F7CnavYnPrb/L7G9j
7Gn51imZ5IRhgsVf/VFuWXrL0lroEwK+/I6mS78QguPxOCXBHAcrtbUw01SCGTaK1vfX3GrXYF1Y
71sueuLYrkPkE37RUcG9ArA/GQ/KoPUYD2LVhwUIjeI6YFZIz+7mxZHv1JTw+cM5jNh6L2IHdgP6
oTRsYmQ7RsrcgKOv8vNaWZtT5LAc5d1FHXz7dQrS71bFJbf6f/p50U63VT+J3gRbxckgfnwidfdO
Nm+2gZxF3A1OUTjYGYD4ermt05LvB8BVng7vxkwKVpBtfwTgArcc+SFzL1FRqlvuN+804VByEkwE
9fXR+d+zNhiF6XXLWgsv71CVRp3BbZFU4Sshk/Uk6SBG2NpX7b3Ygau8Uft3c+nvJAe9F2NfrThn
utvRGJZJWdC53el5WO2mJdx6rR/e5FllY3EWiCr5si6tDzJJizwRKXYmt9Ks4yOrP4gjynhtggnW
djklo5If/t1UzIIA0g/VPs77//lSaHcX8HOOWIyBeW8iM58e5nrwKH5/6rZ4QYE0DLsUGsFaO8NY
a6Pef0a3pJi8HeXcTXVen5g0eM6NahBWMk0lc9opIpNsXizaS2V53hrElgX5TVc0/C9Cshxe0sZP
jFA4CbvpwKNDNvikQx+ZXWGzppk8wr5vDqX9vNjrFjNHy3dr3Kbz9ArWp+ttAb/DRCDvD2So8qcW
DsoDsPqW550ARPyDKJJmWq0EqhdDcUvTsCNQQObComc8KgaaxeEKDFmA7VRwye9IkFXHgL5W4CDH
3dRJBv8WJcHCmXZ/nNKc4F4KGQZ4b0/BjZl31fq+shogqjwruvKy5WQKEUI+p0IegyFuWQEPi+ug
ylgkJL540k0el4kjPuNPMHWPP23JgGL+yLxbUqKMWJIgQlVfput6cQbSCXyuPYeM/DkKb1FpE8kc
fpx6ofgojUWPwe6mQ/o9AyBkwLiSuaap689ExKstwZB+LpfjmxNBVAuA1/8KPXtZchtpsGZz3UrM
QFLPQD2BGFV3nHI7hcLkT+/dwdUr8xnxI7jpTMJA1zf72VVR3e8bn33xmVTh9u3aP+u28+clrkZd
PHCcJHmgeq6hiqFFK6etU5upBwOvgBlZ2Edrb0mwLU6owtfe63dlo4usM5ogJby7sw2kdWuWcDyc
JM2xbZd3C6MC7P6+3SFHA3UOesZnUye5oIvZbRkO5b/qlZqNTvrIiPzEHjophJAK+fEE8YzxjSCs
C26NOEajXZkHHHrMCEzVlE4SPjK8pnlVFP4ekLlvmNn7om37bbEOaWoF5MDC5wSBX56R8Tl1bY6K
Ld3ubCBw7IZoNQShF1BvZwGRsA0swtwyWdQkwTRRqRwvi7Ii/dUsaxpj0gnH5ayEODwj9S1/JcsJ
zAfwWxi0r7+Y1UKzq7pgHGLgkrO7enulTE3u9Is5wbwzlXQhqa+vcfLWFzDy7ZBop2WPJOgMZjV0
IT9KqJbbpIZQic7CLuX66WviLLreTdLoSDuDsN4Xyn5+n5FN8HFvBYUFH3JVo7MFA5EfTDhvWzlO
WgjuXETeFU0iRvIjbrY6Z6Ww+ov9OHzH/NMhh/wyqDTmidkAXSpXYBtxqwdP2m3mr8nn6KtYXYOE
DOq+ih3LLD+BhRiio3BNpEt0c8NIdP2PsTHM9B/MNKpwtJkpFanzJLqfnERvl/kahyPUgI1VU4dW
2Mn34Jz/2QUWCB4Uq01FabWM+Q+nOYUnSB5L50Z0RWzpn5JBPXME0JXMd/iQs6ATnV4XhOCrzYIc
1waeAqV9DovDkcCc9BjiV/1eUDU31CaXxgQi2lNVCWfpDDpFKlxI5vj3kv6k/EBjA2arsqmXDud3
fxtfO62X1cWBzGmSDHbnwVgkKUDfGP84DMsBvNyzEdWPrCpZuO2jXtF4EdglV8qb6wyu/78NCO6Y
RKeffR41MwpeBZPNy+rnjNOCBu+/5/MCevtHfiKEVA3Dd8ylgWV9dYUrFJlINsvn8lsCNT0TT9PH
2HR41kAMrUyP5HnI7me9xbAmJ6y05W+D+J/Y0+dmL7mCtgsvVcymG3WgvWPm5DXzV35LZ4M6zduo
vDgswl7DqK72GG2qd8Ps+lDA4JytvHTnav2q2MWNwHwCgUXtWzrzJpkVlYCdkq79wur5h1A4vx/H
olfz3IpG3jnnjGyFxBX1hIxeb/nmORKST1/IcnKX2yqfV7We9jRH17eBwcnXAuRrCPKxMn+G3UZK
w6qmesYQuod8GlzwkHeIjdiXAFuymXpFG6Hke6yq1HD8nrKB527kkHo1mxyKhqWUMvtgKCdNZGsD
3YS/bUe6FDiYg56tEQBVi/Mrs7sF+mHxsXD63rk/XN/+11tjlF3o/9yzty+ZHRD6Uh2+P4DwgYhj
zKNbUxshav2ObBuzrxp/xmqU7iu+yF73RhvyBF0+AisW3CX1DQXI7Gkt5XPXrtKZAmwJfcgkVHj9
wDnWfe/Uz1JVQ7aYysFTEFTKXMt7kt+gCK6Wwm/5T7HyBZ2mFd5Ff2QmN8cxnmdQSdikSeuqxul6
1a1cwuUhlt7loJ79MnqilpG0VBqjwRjr2ltKEuBL0rGV542IfA0eszVg1K0YRiter+KlkoBwNEzh
2P1UaR40kZpH6W9xN+cfjZXbF2530Qy4wHz+OapttkJwCNUfowS9dpd1Zd6IyVbngtIO/U5LdV3B
qh7yHe3nH1OLE5z1hfGYuhuDC8vMXk+66zDn7+HNSvYtNw1u4f3bMiwfQvLAcpzuV5aGxP7BeelS
f1QnXvxzLTX6GNfHDUFfGLzzdgmfMZ3RJb+d9VdUYiEViuB82qZ2zzJRWgKTfhfK+KJkBNhabIT0
1iM3PzrDaBHN00VTB/zwvp8fcYu4Hfqtzjgmv71/lNmDqCKwF+IY8zCt6ePH+mVXrnel1VBPJhIJ
buP98PpAxPB5j1G2K2rYiYVN7ce+g8DSaxigWz1CI2CbwzDLiobXjckQsl6JWkVSXAVUhTd2qA5Q
N/MUSIc4R4aJNXcEClQonLVCSWsMgYQRos4w4RXTMBIWVvqlfypIvBLMC3gnXN1AMn58Bkewtg79
I5Fj2+V6+xJM8WpmYRApzdGHqALQqw0tyDA5zHp38qyOkfFwSnwPmdzgQx4B4tg4TM7jjwk9O2Rb
oy69e1R6PoxZvoVPOlCYZBX1zypjZZD6tbkui/gCNN2GH5eHXJqD0GgBJw8LazZdUrcuTV6xgKZR
Gb4AEFZmhiCzRLOc0aRq+srlusflZKqAgOdHrJqdSaA5GE1bNuUAmF1hwkpN8QRp3Z+tLjO1Spcr
3n9Ke91KRUORn//CUI++bnuTKstuuI+kCQskYbXeSoJK7IDiHGOw8Lwf0bSI/Y5DhGTzQ2eaPzUD
o6Xdp0s8hEymGrFRLWl1EftM2dmTWFj1sXRPLkRn9r+JcmmwZWoi+KI76ol6PcdYpH6zXo3EH/3N
DLSBmOWlVO8QADHeFa297GbpDUxwAnPG4P5KaauNfnD6s1lIe2rLhGDuWoUVyOi85FnIBmwkQUY0
k6OXahWUMCVq7xKpcBISyxIiH+NllqIqFIsgWyTPSC3lW0vJLQMKkyzuPT1rLjgZ909ZMRfFrEoe
t/0nTNId+KQs9FPck916YX6Q8mYychsH3GdErtRV15/Mvq3Be8dPo7gy5m8jmcx7gbSpSME1R50j
8GXWwYpqEMdNKkDbM5ylu/e4aKYyzKYeNUpi4KUFae7xqNbUQHGOZRrFVtkGredwrYwLgTJK8u6I
l729APSadkuVxtzTHMCgqui6/g90QuosDlsi4OLzLwBlXfLPMeJKCJ+ykso/8jPMnidaeQr6QF/4
sPUw467sHYW0DZ87iLu6rz/4D+qgBqi6A/ycCPncQ5NQoyAl6iuHPn0/IBkESsgQ4GjOq+tQchHE
lhnsK02P0MOZ2XJHLXXA2gimU2MK6eEex1UPJ9sx1lR4du6yni6PwtH2fR3C8O/GQcKLJJQHkekd
cmlG15SP7LFw0X+gKxwXSMqxWnbUhSwneHku7Wj/V127kH52EGKJKj9WdzRMX9vpkqx3XHH0ixrC
RqMfneSvWNoiFYkrbi8wOeDyqV8e5zGOKNAYa67WvLSz16JeP7JxSex6cDpioV60sH4v8XHHDcp/
kQenS40q3UtogRq9/V+m1K6/YJ6UBxy3xZbn17fk6j7l58zFPMEeQ3F+aiUg0MzEJLX++YvexGtH
ixjEj2ioqt+9atOj00pSrPO8KVE8LkEcI/HFmpKNBUwRl4OY60gRy+UDnIqeMN5QEW1xRAUswcAM
RbCVfGAUOlgpl8Jcu7kJuEBs+n9HXWovVhybm84mBA8UgcYv+pWShBHfK/8PdszzBdgcwZTQn9n/
DA54hUuQLnwnQ81L8dtd1eYDkazzaSUDztIjAuFwy4WYpWXvPKJt2LORmkWtYRxLOFTLRWjq5q6M
P930xnzQ5xt9Pv9Kvq0tflKicC14+BdFEL3JogA0cBVTs34gSZfegrTXBOFO89wiYc+F4tpS6QJ3
Mn4pR/E9KxVfDfKA2rM1R3zdI3Si3OdMnjoY/DZjF+jCQhA252aEYcMI+bceHKbeOLrSO8jzbYXA
z+pGQCo9rehBnCMvfT5/ePqm3BCYsYmdpm8yhy/wsjEgPV2EeQoPXWPydXlM7i0drgSY3jaKqLjX
4L2TnxBvd8HNSGhdG2oEDasyO9R2waPiUuXzO3co0VNX5HWQFiN4GZ8dQKQ8Hen0NWSktRvvb5pm
kZs/gyuQMUz9cXKlexaYbXyVW/FE+EPDALjill1CggzZdhmC5cEQ9bqMwl2NSMa2oNqefg83czvh
5NTWBITMRdymlxfsd7SbKFgc9rd02AeZO/ZzymchhVty+QUGVUtM6haCPLsr/jLZFmsfTVD0U88R
wLduvj2lXpUJT/g2rjg5SVd5aeCIfGtdCGfX+xzSzVyabwE250DbtLCdEs69omK7QeXbwwsKCSTj
SHq/7iEFyAjVmE7nZ5CzEF1rsXxn8HN5o6TAImZN/GZV9LAILrOEUvh+RavNzS3Py7cRPTbZibob
ZmGrpRUfSGQcy/X9hCMZP7+C1JCmRtj4N7jtyug9GtyRCK6xhHN+SJ2jCwzdD4x84xMipQ2sqpGS
8WRElqZKRyp7EtMaqeAyTTk8qwpku/U1DAPnjRoYJCzNpoKoSpBExmXSCSg4xvnlYUXvmfGREkg5
Gexku7Jn6p7pVOqs61nIrekZx5C9QhPBBBQceXoJC0nBUwIrXi0R1D7DTI1NUyeIEEDx3RKdCAfV
ERVnXwtKfHrD2dvZpMOJZjeFmMJ1kqlxm/VUScHktsfqej+aPCl/Z+lFxwyZfnEzRGnJmwyB4wiy
BbE/uQOjS7DRZpfWCHwIRL7pCULcaOm62GZzwJww+Sv7pFu8n58Ih5oJA8bae8YXjVdXlR/pZOl9
ESx7O3H+xatGR0I0R5R5uDpcqVRh+FogoBwXm+tJQHdKng4vpmjBbijSwWROQ4/3CzZ5T2xmor6a
Vvod3v7wIpLyorPyIyA0cC5APmbHT9BaH/XfhYeNEoRPgJhFy3m6B9+4czDLMjB0bXLEDs6oIlwj
uIc3zeImVh2tZyKNENZLTpR/Q+5+urSrGUC0yVU4LEqV8ZWiDGFk3NS/pGzJmKq0XwXuMTXBvt0N
Z5M0hO8pp+g4YlCDWEekz1z+9Rv+ofa/ozStR/SmbZQdKCKOMBowuaJtZ128V6+r9uhCgh48ndGb
scwfLimtlcMEJICMZpELrOiwko78bNm0R9nl9K4co36zQe+8uj3ttzZb4QGYz0993jcUVN3393sY
MtdJD0yylFMioUfqjMyRAdmtiAlArvBj75JkS6ApjkpPp3ZlkV/oA0SG7gnLKWUc89CA6cPoAydg
5/2p8FbxdgEtLmwyNvOXtR2p6Lu1nB2HMNMGNJFV39Q1zalpqzcp84XPNT+ldgxjg/PFG6zuBJPN
ULT8yCXZoklGbowI99sFiBcSzFWxgamgmFZqfLYg1pmnNrANSKTO3cB9wJsWXbmrTIk2aHUUb1T9
ol9gH0j1HgXP6h1kEkDocxzXuLeW2nmp+GopLE9hzAzY3gQCUn+uICD1x2yIDGlslKwfCXHq3i7z
SAo3mIJ4z2IoJD+00qlMsZLQKeDXMEFtZu54RMkWQkC6pwf5DLion1hJezzJsKdZormTmWXpGOKJ
NCpvzplXSZSZoeoMI2s9FK4lz+juRx0IDPWmTWfYcRpLXUMB5icaBScn+Ofx6hM52krIDxQZj5tm
hZ1gt0c4U1XSWE/LyPjdRWaGJTF1LeFAq0RIFxI19hXB85EmE1c2MskfXVKYdG0YAsW2iawgUBgR
yAb36PGEpr3q+YjBxKfboFQjy8GOI8p5jZfG1gVa7dXVpR4NCKqabc+FDyDT0kdB/C59/B8DWqSi
xHiTtrstFuSXwnOCrZQxM+H5UAwjKM5m0pdgVZoEYG8yYWt6A8Fy5OknVzfKWK8xu23xQx2QtTj0
tMuEEra73Qwu7wESZ/jnEz+qhQ/uJJPh5Ln6WSd+1L8nmfQjcJoe58tGaUemMGR1ihCPAxCq34zZ
+XwoVra2t2HeirbYbVy+q7dtkwHtC9ZUHmDvvhRB6IbcmDDatA+u/2PFHJ07Y3Pr2OJsdsQrMncD
gv75XOcCHz+pY6Jq8ayuce6N0Xxsab64WOadjqZZa+3PQO5ygr7HvISX52DnsMzOYC7Wp/OBDDbm
e9ghr1RRvoglN9G0ERrJSBamaj0lIWXuI1LtV5t1z/BqJumZVhm6D/PkyzUCgsnnGdkAtG6uz4Gu
abStVkFhU29AX+rip2Nsa7nX+lx313ER0bqzMtsVW7/W+HfSYVE+LmqRQr+BS9JuMxoeQHMmnhdu
dKSqSYFmfdQdx2pxv8MHvBENOFOoTA2AGXWY43J8Utp2P6G1lSeGwCp//vCCGbVpyablwv4dzhR3
q3QBkT4j1HRy51HKo1i8YUlLWcJmdW6Uo8KsDbBSMv8VXdXuHO7ZFoRGchAfyQpwblVTdiXCi9Fc
z92nmcgylN05qaxJgOj9WKn7dtd6EpSp0EcPPO0BpJnpXGPXwHpoEX+eR6a1a+nxs566fayUHQDo
dQH9WoQKpJzdWKEe9zi8gCp0A5AK3Rar41iBKShKMe3Y7YDF2XGpuoE5Yesh79nj1ZNRNYXemRpY
UZYkFaWHZ1JEoeIYY6t5jUJAajd+CQBwrLx6Z0fX14psQe/YqIN4FTmPqCepGJeX7CuTbgM0NYqS
JJPTpWRBq79FJSqpjPlkGuODJMvvn6Iwh2dN/xBao8Rf6ZdkEfoLn/DE6T+5FDZZWG2BYD2FpZ+k
lYhHF5oigqgdcdQg8LfOwcRaq8aSDC+LqSUYV+232PNiiKX2PmMsrJuG+/d/trz82J5KeWE8ASyA
VcjfIwmGhz6GaT/J9D829FbsL/h4pNl5cf1ozjaLtDd8CO2BZZvJQbmYyEjAH1k18q7q5hSvwAFV
LiX9zWoH9hEsylntycKTknf+CZwnfK1tPu3jkO26fdC8uwVBDS2YGJsA/iHFVsQ6mt4TxBbsOD0X
Kj3VFsT2nRtK0UX0mOvhA1v2SG+dg+kA63oMa/go1Qa7d/v9OLPw8x/COkmAoFQSgRCCQU73iQ3R
yXK0rPv/TKKtsU4tK+Q7g6qp6vPYIKXrMPOdEVZZXpbE0wUobsolOoVW8+HPCPfIu4F4YgOe5MeS
K0YYbLBkOjrPMKa+trJ6Mnpn6q76LmdZv0bLeUnF5uEHN8FDXNHqlBn9ggVgifMXP0nY+80b+u83
IDF3aKL+2QTqX+RO0jKPDE73xgbhDSgAaFwNT13PrP96nEZk8wxfFgT4TjFkLpK9/eaJtfkNWMQQ
Jb2i4wqAkB5FmzozFHET5hX4eUvS817jTVHxA75Ox1sKmDRS5Vv1hSlXgQZ7K0DGrVTTrTQiTsz3
jU2AFNiGwMJ4zhh6rw6ShGZpm+UegP06o6OT6Is0zXW6gGD6r8mu6XX8kWEm6uVbxpUiWvnGOLpx
f2kw9lGFKanHwjSwYHws4IVFdaSsoRv8JGj0H2oicKawYkJzwTVSI0ciO1rG47UoO/0hY0DaqbHE
EGlUw9HsyLv0GgxAfWlqkprhCg40Ysisqtt6Ix8pW5jNJ+k+qJV8Uw6/ThA1itRbi8r3+BACeHov
Ju6dP+NJUjO7Vbx6QZ9+OOSVvvDxYfLJFUmJIHhRb1kbzrOE9wV0WOYb7e54z/qdpp5tkPxcftRa
asoT8wDGVXNfI+Qulz1uOM8ULutdAIXUlEYtAES33dctLAbP1LUJ99cHTXi34vf8jM9PhbqAdekj
bAyw16nwH6ua/J3afZVy9elsGdyU40IlpqTujLTonD21ZmGrjFE5A0IApF3l72HoHEGisTwCV5cA
HkeTq4FMUFAJZv7ZTnU6VHKfWAOI0QZE+A8oHJ7ILsGI+2iERYZuj50o1151H+N7gQKoeSjr+M9v
aODtcyvTRUu1wor8EmyNJqnKbZCtaxX/IBLckFTgUD9IfqfYH1StvillK4ObmRBjF3l0+vf/xJxh
Im7zMSUyAkIVY0z+ip+qaBrgWoWjBkA8wPf9L+WnYO/CqKwNnYo+rbY06NgBCS8NbD/Rl0oWsGXo
ffpw7NTqr5DVRxdhW52v/U72nl4bZX1mdUyZ5OilFAMExAgCgmj4D7QRjmRxg+Y+A4oPvqaDj0fv
6Mofcm0dWrtVnEEUQHRjtodlbA2gghBnVN6DrQb6NGhUBfZ/XAPaqViu5/DjdnIwxFshobCu9Q+9
hiRwUIoDZPOyaxzqd5KkXa9A/tZczQfBhOqI/Xco+HfBQz1q1AZDDCU0d6BxaDEL9Vz34YuzMYQu
PNHMa+Mj5dwntIMVxycEGir5WP9849YNGS3Rbz7Ypm38VDV4xCL5AuJ0GhlkuRaiviq0T1T8rhOX
cbtc5sTAwi/eFeO33bifm9/X5bkAn2wW4n/xrfmVHfFV07tJ3pv3Lud3JVloxOKNohfihoYzgwva
Dg+FtEiGQ4l8eTddEbE/DaA8PU71a27zYIBmheTmoJia4Cv7wF2V7IzjLMgi4NQLRFQGIBPlBH/u
LN9aNJ+HqNS7KhqWgKH+Gl8yhJpgxFiqRBTn6UZN/GMAVUrFkeHe46tozcVkNmKDkCaTbawlx2w7
1+NFdv7tdFqf82BK+zYcTsD4cfHrPjvnBNuquEPeONdNYaKZxgaacJl8BeZgG8KP9dfA9l6fhGUA
BXB+XKvVhvVDvpLdmap5Cxig4E8veeE3xXxVcguvhZGHRV52sbyfC6zp36bnbnu04Mo02ogC+F03
2R0vBxTNQXzBDW9hAHQCx9blySZLlijTZwLn3TTWw5bIgYWKTdbTk5dHS3WpdnYR2E6f380zuZB/
lJoWeOOf4nwgEL3u1vk7QNoftKAb9Vlo57xbO0HxxIjut2MqIhEGH2DXCdgLs3UqUIQa0ilHA6ZS
NXwRlpRJX6IT2mcoa9UoRaatrEl8qqKH3JtcZkmN5pvX58L/PDNncEjZSqGDHdOavxIDM+Ro3d8m
LZK2Fniu+xrp6RNkbaRHr5aW9LKT+HSKOapnZGxwOY2Y9s8kRcfg3rCUY/aWFSF6fsRXxQytkyvC
P2hlOgkfW8AmObfsX9ZGj/OGlmhsgqw3xW15YykPh7KjacmNwRfgdj9aFEdPVGYSp6s9+2PSh3ee
708VGAy90xG2zw+X2NQMlv5rh2FCtuldAcUYAe5Lv5IeKu4rtzPt+5GIrCk9IqCfIJ9tvUvKvmll
wux2NYry0oa+cyxVEHDFOlaB+kcc8Et2nXjCWNpap3B1+R0JZnOjLM8yqt60Irld4tTazSh5Ieho
NINno+bntx7vOlx6JpJudLve4zT34GfBq6xMlzvYDzy+wvtTrrqo0WXi3rNqkVHKvDMaER39eTSj
jftxkdWMSi+QBKo9/S+TLRE4aHh9BGAAvmC1P1vIfOUVgNzqrbNw7egU4hvWLx9PKmVVcvHKl7mo
8TFUTuqEGKkySpPS1OQ2bwSR9sLsq7tTDTzwVnwo1jg/yPBq/S47Hc9IW37hjgsLMLFC587bJ27+
C0JDoxfMlDuSOsYH+9UmgKqSrZiN7BgOOrFCvD/hmw6wSAIM48Rhx3ADP57qCy9pIvmCf+/YrVBX
GpOHDEtVp9Y+InDLqnUWfGaewH//j91oFxsF8I99fNzoN7oDBxBMBxKXvW3twY9sliCfuXArWdGf
B97znZCN6ieRLxiFbHGrzghMh73yRvXVlbSft2fn7tDhZrNsfV5yDuivPNnIO297pamYc+6RGHei
gaxzyKR545lCo3VusJxEvA37sVS5Lit0ghBghp9+UaF0Fl3FLz8dpy2y+HY1F5FP2deFntr0PApX
lwTZLSboOzH125n/m4Xs0SOVHVkaUVUX1+5OfMDFiIxy7gC052eAKKsfxkib55vM1s6Vh+zGP4o2
lKc35LA8cMbmbHLhzCJFh5cUj4pw5giUvlygXExhTARONAHfKzehy8FucZQBossIg9+NoleNKHet
5cyN8wEBnJ5w/jZAKjXYyUyAExlVuejDKbAiGg0E4rrn5+lYwN8OxsDW8ARBIkXOuzuZr1ZVHL5k
CgeCWGFxicDBxuTWMyibI9FpOjvGqQBWAllrx+Az35t0EI8N08U544x7fxcxc35aVNWLxS+1onG1
omRU3d0AF7LlyzzbDkOhtEZ55o5BJ04gybudE8vZV73mj+bf7wkvypKWoN7UWp7IA1jXG3u00GhX
5jGtd7nSSxYcOQ2k5AwxBbbDgzuFXQHKkHuvhsZoGO1UODIsssnYoHF/mK3OaK6qUh6fK3rUFeOR
lXkuXkxsEBjPlRkEXqYy5zWpmV3i6sEtnHWMhH50FmHqjHdyLEHIlWLvpDtCqemp/Jg/Yb6VAXM0
MJ0XWaVvFb4m/DeDwYU0xIOdDZzH4iqZLQNQussel8jPhEOCYTssxtyaikXT6SERObRNykDEinhq
F2A6aTxzBCsFaQChDXr/dJgKrMvr3x6BhDPeIduR2PH2WnN9fAItRxZxZpsLLgeEzXVNvrob0D0N
MWMgBDwFXF2bihwONd0viJ28BCchfyTG0WcE2UYNWOvGTdZVp1G6NT5O5k/uV7UesHyr7zHjyQQH
XD53+20773DVw3tft/JT+Ls5SqRdOdvCMKrUmBolp6TWaRaqu9HiJXJcEtQUNT2j//xa3eZYy9TH
MlESZ3Uq2Q/I3Vj9QlReyuaix9hAPGbYD2NPFmTuRU5urYuLj2PUrDHLDug3yx5XbN6g+LWmsj2S
GYPzYstbW/dVvo2DhBxFJ1usvroxc0c0bzvPtI1oIuF7MjxOER2pdUAMUCn3kkTTXag6v0nZ4FRA
hy1YiOnVPaBYMQYs08nXgWWToy9ikKNiSRmSBaF27IcnCGoX+pnFmEh2kQUWtypLxuYKgkMwlSY0
s+oxHm8R9t57LT+Es1uUqUIzxpVfka6aaFIUim0wLYAtRi3lAJcZ78mzDTZoTSbil7Jf9u4vLENx
+oGfyhrH8a7Q9VCyLavAvJphAEpk35rXldJn/l0oII28YLPFmZ2LeuSkB2+2VuQQ/DtYcp64LLao
rgxeG4GpZRLJV1w6VnFMGIyDDWj6sysPeIBFJGAxeiCsBfzq2bukmZ83KuLzIYNET9UMljE+5gMO
57smloj7euGIxFWIZ5nt9Q5UF/HF01WzmltevfLxCJOs728Frt8R/NC7yAJgWI95pgkoQgebnn6f
TMgvlHIRlVQsQiZjxt04he2SDascNbw/PHsw23N4E01Tb+zC/lxNoBl1MNJKbf5oy8e18bqlO69F
fRhsr/K2AdbodEAzcm9e98j8uPT95v5eVHX/JNJ+JTtpQ1IwDYhb1HIrNIfpTwuEK/3Rb2aWNwKp
xp/tyDI+edLGx5sf1Gfzzx4YJ3lNbLmar1+N54qmxuUXPNN3yYAGWzFuvR8xjVYOJCGJsX1zo21N
ZC0+7h7tai/VECcAJso8mKiI/pQhFRFxuDNSWVVnh0TKB5QwkYBMUJMJsqVUK1ZKoCFCG3/MnwPE
eBv+GGG9cUmWOgf6wPvSS6Z0/VMWiB+bsc1wkv5RU6L08XevHWOjOv2oFRw/BfRUGgZJz1bwUk44
fYGCBDtlunXIMYTZ/Haz6WdpkVjFX0YNXCKYKzSuiq73xAYqMEqzqvc4Nyo0TU3mWjwmJJbhN483
SktwCouD2lRbKksjCTDrHqy7hYr7IONMjFvT6IDKPXZzk1pqOTyzEy+dBDzFBSCY2GS56MwJz5pp
NdapcOm9wBtBXyoraD6quM5B8swT2B8nZyodmQDd8yFcccfRyECuS8IdUIDaElrRDP6C6Blm8Ol+
pFjNvWVD7oWNNbfytk0s2FZ3b1desGNuTDUQ2bV3xtjP+Kk9nPj8L/zGYlTJpx/Dn3U7UAXpeRaG
fqCyp4XwM2uL3KpRT7MkTGgWP+YH/rL8nYVkTgQtGI+d5lyOLWsYI9pT209xuEUVfi6ZI4YMiyQT
oBDd72ON7ENS3tAW/XjhR6buNKQOntivfpTuxLUdj4VxmIr13ICW7J/+e0Esf2YGBgysTgpBN4Cu
XJM1yPi1hxjrY5WbwXiQrrNSXzXfdBLXrjHf1vRK45nPcCLW/FaDaz7TFnoNfNkeiOs33XCJzwxf
D8d0G5SjlXhmquz9RSRq3av7NjNc3dyHYrtt23/Dzmo0mXVHb/EjjEZQ3RP3D8GtyD+u3/3EchVD
Zun4zGjddUuPNfx4I5xeeWaccHXbLmAskAthM0FWlqE3KClTkzra5iFBNf0OixiIgZE5hxwYG5Fq
NqGwdSjy0kGAhKjvXZMyhzNaHzmWVYolzKSZc5DszGJoZzxx50agsDN0j1/31fg5/OEtJ32V5b9s
LD6nc8vtTX1mGZsYvxQuvNK6fneRbHHOVjnnnXwigEPvF1GvvDpHc3AkOdImYhMMcFLUxrIA3wVp
J3iexcipJ6mwWBaCc5YrD5cOpquBAYeZMijm5zLLuh/ChMRTHyUSsWHv1bEfqn69cVbXKIuNXIin
B243LODALLZ5l6eW5Lfha0WGUfEuUJo7tBgQoGfGxTDBAc/UoM2ONF9ywRCM6hQfWmq9ysnaN9UM
UZayaWDuajWShlIm5+O3zrchW01uuGRAsxf3ApVxRwtDt/JIouga5wBU8gXe9NlWRidSd1GAsDJP
+y1RhKhqempFtaW5fdnOKb4DyvmaUWtkEhXLxp8oDlSuVfDKXL7iHyaM4bO/J0d+DRfoE3ccT93r
KbpG3CmjZiyfa9i0J/fzYbigFsKfGMkLWzfzcDY4Z7kU9awEDluTMUVbC4QWDZ9ejoW7ty7k7lhh
Iys4YdIXY4pCbwdDjn+N+rkJTICjPrDsfspgCV1/TLWtYjyBmgBNeiSV0slMKXk3WSgLR1W4jvB6
aVSXFIrAkWJhYF6n6tVnw1bdEaK5W/X45NDXLkw5I6S0hQ2fwfRyXkmnlmq+lQgkmezLeOVVVPk7
7EPlNx37pvXRgw57EOUnAIMC8XTp+DEJ5SfIiY5rdUilzOzLJ2ab249jdbyNPu6UVTrnMwXCtIzP
yhPI6ORmcrgJH4G6Y4s1/eVocR8NDXXMUB7qczhmoYK7vyeA05qjEyATobI5Pc91sgPdco4PaAkc
YAWsotRM8+ISd7BzjZNAZSe90nBpSvOsYVHdFRh8qqCqAHlJxuh5Uki+jaqQ9TkFb3mIBgPd9RX5
Jr/lR0TC8ScnWH1JLvjo8YUDKrRCZ5J4tuTKBsj79Vwmx57AX3Ie5gICzrAWk0QpTOd76dchP7kf
yhb0+lj1W6nUCKHOhsXKWCLafDAH9G4LFX0KAXPAsj8npggM7YU3nMl1dfTqdbYNO1Z04tu/4Qnr
9OwBAnaTopCAPvXdRQPsuI9FB5iMZwQ4HuDm0emjsOka0mdoxXBDxngGALM0YFKAmz4kmke1ZTup
zF4k2aZ8UC2zE0b6J2/EavUGCbrQv4vS3pgJt2YIXSbi6BCKilVp+S8j4jXIENc3N1SkBoV6yZER
tIV5l7y0ikKNRiYMJjTPJ6ghUrOh7zGoO1HsumKDXgvXhe9pS58ikkOqS4DfNWJ03ijt1lat2GPm
cc/7xXL1+C3qwzJvCoagl9Y1pbVcL95v4Sb/D+yDeHfe/3PXio27P1hRi2aWeJIlB6wAhvWSjJ+6
8EH+weu9HqElSvJs4lwQQjdcoHVV5V5QMkoqrXCO5aYnaWX37HXQOtAwIvr2jQPS/acasxGoeOyY
1XcGHTmDcLZ5ZR60VZCOFK2zBk8qpGno3ofEl4rZxMZs3wnJgbsWhYnwHIp8C6lk4ubUx2CPotiG
BZhE6GGsiGAl4c5ceIUg2bmE4x+qlOYP79zXLzG2Jd/iI32LLzJvxDJBIbRFq275FAPo8faSRzS7
PaVgmgaKfv2zU7P10JqInXJtzz0PV7ym0IGDVdysh+c5Ki+1JpszUvJQTouZ9TfVA2qBOn9Hqltn
2h6OysQKDfq+wYrfycjWExkQvUudSSq9nW7X+Pw+4IUoZl8ssdaCXLSWKQ7Wkg9TBfhDn/iouwwl
ZHfAwWHTXlJkfhChKcRnVnm9VNFAN3pmOr45u0ZyPlZde1yY4QqNEvPKqMKgeIbffNS0UPDHI1f+
pGimykKqvaiMgagbydjMYVI4Iiwy7zxBjbO1Jb9VIXlhazRg+ltH/sKD6bOO+1HyZyiYw3Sj/TZC
AOeexW6LNr8Y/cnNce78mhWw4FXty2NjYYI9lqLn4fz97DaqJE/oojP3eBH2xvDtCv5DOkJCSVxC
ZuLBxWewt9UZuv03+JnqFPaJ4Yb5X9tObLcjQV2+/+8FaWndaafYpzaEU3QbmNbsWVMYqLxqS3qJ
lCJ/LoJU85ZKlth//gjz3Uu0lju0zeejqKOZ1powQRl8VcHL6ZgidKuJE0xMrVl1c0YDxRcDEUzZ
CJNjnVTDZnhoADgww06kH2g6E874ItrULmzszJ94MYb/ll8U+AF8S8Q8OEgZpBGskztBbSQmvAx9
LLd1hilYXSRbKY+UP/SUxhCR3feBEcPObywiR3ztCD6awpb081QWZ8rqCzCg8KxDgNRxXW+5NSTM
dfJaauGqofjM02AudFrDoxWBDHJMTW6zeL9cGnAz8o0Zfh6R4ek+VCuCcdqH6UfA8F8kFO/FRy87
Jdm3DjeEBKLSNgtiYK7TqirLTRIImSNO88HBEo+nIcRtXEV8lOx1u3esXEx2e54Y4R5jlwBUFAO8
O92IIbZPytmxesLD8m8ZDrr3sVmyxmt8B1r2NKn7gZahGzEDDGihY+TBE5cePV3mOPYGX9hN0/Qe
0RR7xBA9MgLXeBSBAcIMakVQXFRpxcSmCSwETBdVUiE4aIUr/Y7WQVpJiaiaLdRnkXOcE7zMfo5u
4ErNJLkfrjjCeOniovVidFxVeX1qZ9gAudsMZgpu7JLnMSTqNFmBMHF54hf7EklDkjNcRkgLnyV4
EV77Cip4aZ9g6yFBuIOEy6bD5cGKbH2plMkKcgWvo9wZaxG974yKqKThhqiKeqW7+4xYGgTpnbvB
pMW5yRGI6mGZIXuEMmr3NCyCxvRdsJabohTkBvxKQp2GnKe2oJNhad8rkdbqMrWE4Y3o7d+lFUkB
vD308ueLj+nMMYuFuFQulG8VT9Vfq05YrOClntTkT0Dt6N5gjacK6rjQUtwpKdwu5FHWMONMd3U4
jZBSleFcsGmX9ak86ylB22uN9fdSpG1iljIGAuGZAURsNMtsBQSDqZ9vbpiBuUH43Ux7guegkAr6
ktvybGrZDbKS17nHhNYB8nJuXWgTXb36by0Ndw1+aS+NmRw7blg4HHSTwQ2VPpcViPF2ZYq+wpNr
O+n5CW1t/ezulrVxmLc6M7OgYXqSKsZ/sd5fzasMBVIle1x17xSACHccfSu5Te1o3OJ0RxTR4QvV
D6ffcseFqRZaQyANrSde8KGRkNkzCIegWs111v0YqXc7ujx2QWL8mB4cd+cOmCZVzlwwZ5TwLfCO
Ob/ty3A2E+ZQurBnklAr8XKO48/H4HNw/GMpIyi+yPeYHQxqFxVcVEDKqSw9bg1Eel0Vw/k/jge+
3DNyv6ur1hZ4fHbHdz7eUQmPVswtal7tYPt+7UBKaFugulhevLiQlbEJyyiXAe8QTnlvJoKsQSA/
OVq/V6LjkQS6HBFMtovyHfx4kqIRoBWng2uBIkJ7vWWMbCu/1rk8ecvkabN+2eu1l5u2V+Q4QJCE
15Fpg3p8JIvRPd/Ew/oUxI4ENUueBdssQXGPEgwYz7c6abnf6/vUIsAgEakAru22dJJzzoTC6U6+
hJ/iARjTRksazEAvWvuGBcKuEJxUdbPhAtd3B0apDmMgLnORbafyKOgJAl5l/CuiNpGBJliJDfD/
2QiuZyMgTRigmfrm1hxQH5ESsYxA6fDsaDHw6vIUmGsXUoQ4FzBxgAWy8d+b93nGI6fvU1Q+EVYL
nd0h6+dW6qeTLkTAosy+Bg1PrijLB7+IbaEma2M02py53X7cts44LByNGjqKjXS2Ib+PCyE0YVxU
plx5wAosxVKhUubDUnK4+0QznjzqgxFyuf6g6BrrC2tzj+KG13vDQoDiw+/mU9g+ZrSDkQR02evH
e9zqNsXZx0VK1tR5uZ4kBOHyLOxPyU3n3i0tY2VLD3Ey6x3CjO6EDBVZ2f+157lbHpn0rOriVZlB
xDdwIYYrgXthcGRIyqhlhCqDaeAyca1xtmQI/cS5ZAxLoTnA7sgr8fT8tRkupKgti2jAIq6awHuB
43lEJqGhuX8lfjnEpzso9DOKfsaRg2wN4alMyhNRrbMDk1VsyK7HOGwoFs2Adgh1b7hBaH7ktfJY
z13LHjsle5iPnurG6pX9YvIZTEC/GpyrX+KqE7IYnhT/N4PGMiRW56kB1CqDhExbeH7v0LvXEjLp
XggKb6oDVy/P6u7RI5W2SJ4NS9EjynOqWivDFhplAOiKRtqTPj05xvZnSP+dZuwFVKg4h9SsuN7K
Ma9hQbPkZzh2jNuP5bVgPD2dPHjzpM3ZijBloseVPHQ4RbawS3zek273raQ5QjEN0STqHGEB7W0y
n7Mj4SuXje3N6Jr5+bgWnoU091xalVfxScKMOSPClhUO61Yqrq/xLfqxRzRG7QgOmKyGDPRF1uzf
OAMKJbPJKpwpaNy6AOl++Om12wPT60kV+Ztij2m5g1ujY4Z17wBlCbKDHc7CJ3lV4dlr+i1pkY/z
vOZVC+OvA2j2bftQEredfL+YHJgKWdplOcaOJRZ4lbvVd2iaTutolyRIO3JSQAVnECn0bDla9mGR
in1z5nPkMSNJn8b87nh4IPEljxa+rCqREyo1zhYM4MRizkFqo+NnbOE1L87nrhEIs6E/KF8SbTxT
uiOotU9+ntcBKz+FeDT7MzQeH5dTOQvb6PGxm2mKnxLdJjNnzfTie0GadWhXVKwaM3QcKI72bOc8
0rObfSbp7H71DWOLn/vkRjdN9z1BM3INRV5SwjVi7Ms+LLQ7Sj4EoxqaeFbcJMBn2+x+/uunq+Qc
mu1mwGp3cVBA971bwq12UxpfMrHpMFswCbbTROLG8IyxONsOE2CyvQuqonGszVp75dtUHXwHb7Xn
lXu88h2HlNdHaul8Bq1j3tATHXI2v3sC9RqySAQlKdQZ2hm35wn9kidiXiOgIrHsE8nSABrEBFVN
w9L26969JHDKwJitgLQbyFzkl7C94Jyvc5XDi0mJMENPxD+c/WeBibY9Co6IVG2dckcNj3xPXMYd
hTdwnfSc3G6u70dXRcJ61Q6Y7MlzPGq8AYHq31ojgpCVjcM4+SMcG3wkFr76izbB2Nre7Ro2iCjR
0OZj9Gzgm/+GtOT76BjpfpnIVLa9THfIMfpLMr7PYe69pb1r3J1ylOVboYLKr7awB5pwzXZ3aoc+
WA2i9Yt3oHyZFUiKb7ygcKEuJn4lf2H+P07VfqhFYxfgktSCuQgm4txjM42njPczUs44AK1O6dDc
g5XChtDvm405B8usibYIfpfxOkqB1z1tSLf+OQF4B6bs+/UZ2NepjK4DCBlj7JkKxOaK9UqMPPUG
zW3cGkV7bemT0pGDHfp7zOXGBxB675S628J5rVLeUYmXXu34IcYIgPFFcVGdtV5FCpCr/5wKFNKL
qfL6MdP3D3n8z3nffHS/DywrxSi+Va7lwR4VDsOx8d6ZBvx7kJJ8jmdYL6OD1QylDh+zsHE/Lhk5
WE4aaF+15qAudoYqUxAlurAwCUn64DlouxFwV43XOTQc3hIRFqDhXZUxBDTnQ7tpfW0hewBt+KXW
/3ynVmjT/bFIIt7aQ55EdmyFxc+ts0UTufgsYEsj9qF83YX/bFKb0DeU7neEbvKqaF7JIdjzv7Q0
HeOqin88u/xr0rQkB4j9D2hOlbuwgle2FPerupQwv9X9G94usCOuNnY8vLAwAvixinNIHyd/rhzL
41OUKscxigM5Di6ZpkgZDaRTVGePQD4yaaO2ZxvKDVEbxstnjRrQTB7u98teZHx/dJkE7tgfaDEB
vtzTtsMP5BZmS6Q9de4YFk4KZV5SsRGa+s/TARAmbTnM2Sgfz6Y4RFLIK4qV3DcQIOpS4BXRYgXJ
mrDF7g7KTsTUH5rZLs29T8q/7JcSqkV2U0CSv0ENE3C2MXscSiUkc82bWepNXwhHmjhV2+1QDeQE
i8YwFeD6VdGqPTf4vMM8C9LP1LX8PO9WDWgn2/bwEtBQo2kZae1TAdYbSSPHrpgb2yn1vDMUJgf+
qQQVSzl0J/Nmlef9ZxamHYDNA/jfS1bWb88Mphdt3PDAmR+i8vJ7ldjftW5YOid4x57qfgTLT2Rw
yp6hJP+N8AQ3hYOPFXCu+4SBX9ENux9fQm1gIdoKWBQH+4Mpmwzw9+uzY/xeTq8530ATUu6fgW9+
abn9/Hg6a4wA42Ne3PQu6KESu3teBzZ1zwWXnOHHqoruj/vF8PnK6+pTVY+WZ5sBqQXjSvN+MwWm
HZan5cXrbwmN6YFJfvJl2rwjquLJ1zuvpn18Wt3cFguUpy5VZFRdoEBhCZQBvDkD+WGDERTCAH3v
P0pEqpQ8hOfZZTy9awOWXYvvNC8E4761tantPA6Qh27u9k2mNhdIjnzg1EdQZ6CRsEKdwy/9QxcX
yYhOboYU7Yj1rEOF0kGxMO1GdBv84Ta0yo8fNIsX+qGIV7CiV//Bc8naledGXcrVbBXtQ21Pr98X
aTRmpF25GLzOjd3MmsfisYmj+sQj4JWdiN5jQM6EzdPTNu2UoKsPA9GQFjkrvX0k/LGBGdS4eCkR
bVnAFPKvEPfrh98Cj1jTGHZOwMMipeg+xKrNvrZOreBMHyCf8hFUMnJkV1fNG1V93A7aXvJTwbpe
3lIUwv/gf1kdyLko0HXE5FjQSGXxo5X+Ag+ohwJSmJUWnUuz2ldSM3GQURv/wqlnWFYd3eICQ+M7
49wvExup+wCbz8vxbOIhmIpFkI2Z8ODaO1CLIu0pwEVYYwhxO+LhEC2d328SQM3FMH/K+r5gvxp2
ro3zOvNag6Q+CI6PqGRZ9CopsbUSK6F+PMYa9j5ewOrbVpnPYn2lbrFfWO3u+cOuMVbq6WVM5wvn
8iRVZVX501ZCBSs2jw3s+qTrS3sn3fJwlKl22FnHrEulkvgtmkAsO0C3ndh53T0dMjh2Td2/6Hve
4opqiQ8x7k9m2IXdXtPYrSd2FO0gKfjJtIIpNRHHj8RMU+vmCOpKNGc/Jjas82p8pOZammL+kkHO
4aFQRVAeu6o13bg38nHoYVkKeLQBu78cdpNKV01P+6FPHWdjit4MeTcArsQphULc2MEjOj7j8vQK
5zLRdmzZAnzuzfiEenZx4cdLyOypcwHDDMnAMN/SMszVo6/UDPPsrGyoN8cs0OlumVgc9k6fPeLI
wL9dZKGxcksqohYRYLUmwHTkOdBcr+ZxXmIpFZLAjeK3x+6EIj9ZQakNm57h9EgtKR/PiUBndLnd
cD73a2UiM98N9RITOYqiwe/S7WbaI6G9vC/TNLknAyHG1oVg5vIoY+Wo93frtkxO8ZVpNZvjeWXq
nXQXHPEk0PQ4R6FnE8txUc2FFqY5e+oF98SE7wnyCtLnhesxuHBkYSfwPAPIDAhRm1ZMGNScMvpq
CYPljpp3xmpQOIwpCeXrK7TCFB7UcA52rXV5LNJMPMzPpua/P9lL9iIwFrQJCwBaq/TH2k2ShKk0
4+2QW5uo1ME/14rETVLj+hQHRGQGwnfic7sI8iED3XegeFxyn4m5seNxbAqe1TcS3WzkxQ2DWJ9j
93XrE2d0H1epsT52UJKnHjwFmy5JSZlqzXdaVrwFFAHsB8D9k+epAGGGmTk2OPEWgTPLhkbEIoEi
qMbD1PRYVQC8su1SpbWb0iBnzztH0kbiWpxbeaEyZI+0IYmsMcw3Ml5zJ5Q4TlxJiT4F/mvFGeMH
+THkWaeBh0h37I27ZlyVcMW92bFcMZzmE8QJbieP5kbJlRO3JM22FZJ3XEjLhsovNsrGF2e7n7wI
4sB0cj3rq9ZQegz7py6OwLI0Vr/XPWcYroE85QpuJ73/ukWrggIyIziu7LXaNccEGUCzTRtFrTE0
7OnYLwTzcC/5J3qioHs3y2zDD6R/8iVCXXpKVdrms+bR66VjaOZ3m6VkgFX80c3m0E3aYuNc1Iab
7tMIdftORm84/F4GHdBTUZoORxEj4PFPE8MK+HUeeFG1pfeblaSfPnFHmICzRjThJg/liuzEZO4c
dQOF64CUNPQdJy1MfbCGm1wZQrDa6TVfWuNINdwBrIsO4VGH/izpaFxfMv3G+H/s8Pn6TH8kxvR2
Gg1izPpY3jZ62gVtezAqm/9DHt/0RnKlSHjcA0KCDgN6T9PsgxFvAVelsaX4FUIwbWWlg6vYm8mZ
T3BcV3TN/ARmTGddjJ8sYu5oV9cLGgOcW7UsWF3RXEhhj376bKxH0uniraSkhXVkMi94+PKIhO3E
OCvdezi+1w0SAZTtesAlnABdCvxpJ7RjEYxGnwIn6ICrcOPFiVjYjtg6c3n07deb9NvWAUKdCm6w
1/J9KqKRKXgvNow25KUzUAY1bLs0AKjt2fErHkN/BvvevwfGvB5s/1THCEFl46FYIq4EK5d0IlYm
RvVRGUqlvswDkmJNzfex3fmCv7stITFaMzm6Qpg0CjRTeovERWKL+XKkTbkDaqXeXVE7F6srGwZ+
nphHR1M1oKEX59NE/zAdSasea4Y/xV9zggVJkJbHujfEXfB0toQvkAUUZQMR9BbolrXIdo3mNfI0
6AGZca52XBAA7pffu73f7eqgkWQZDLKRDbqooxtkXFmd8Z9J+cNQVVSebdYSBpT5jp39AQCtkuoO
oerjqSWP1L3JsEdnJcw4t3PekuKqYnLqv18vW7isC7297JaafC36ZZhjFWYgYV8LYInYqGANa6BC
+zIIR0K7PqE3l9RpJiHfAL+kAo0VPt+63G3L0KP0Cnqb6CGYW46FQI1UERkZrmEP3M+DwRYkLnpk
OdcYcSa0fmNj7If7srrShGVh/29+rrzyK/UtUPLXYLoFL7Gt34YnKR9vHcFP/TBbJAumJoIwy3sE
1D52Foccl71jokpubJtakK+p5nF/67TmpGTWnCHSR0OM+hjisatlRpakrncOTP7B09VJbCKII3ad
v+JNzi4J1ne5jiXTuEZv1D0Dkp2641WhIRwlJKrw6vzOs2IrxCXwCNUU04UNTJco61e457M7SJxo
XSDWbEEdyZu87Jts+tdCzXzv9sAFaZ5x5rrgevNeI4LinCMiSW/VMujkDweFxBhZ/ct5n3nQpNya
5938CfJlQOL675EA3dv0VDpYQT/uVHaFGbWSeF3kYfc2HUI7fY/kehMaJve2B+cqN/UuOISyze8n
cJ1JIHC7NdFFQl2TY2sYJPBxXcbHHOtvLpcBXMqrC9GIHdS4LtE7GeGcQBOgfrkZJ8Yf1Hxk6Wng
O6KnXsyPXioZvLIm4PDieS4phCJ6l9oiltMIloYbf5c/jLUo+ClUrFrqVOua4snu7OQKoiutVK2V
rT6UHtQug9L5DcF7KiuuhdLQfTO53H2h5g7bCBoABT+yLGLNvCaUDrnWszKOwE/aR9gTWIczxrB1
uC3pIjIE8+H7DrMjA7b0kXbxFQAS2czw88fVac2l4yVJ0x3nvnUjyZRGlDzWEM7wGf8wxjhS4El5
a/0KnRgoo7GlJ4ZtYDfEn/0Ha89Rboka2y04zHGoXAzenFwXg4QAAChLWuJA0WrhS2FrBZMCxsCz
cv2KoppvMuYL2xZJCoMprc2Vu3yvGxtZFCKCgbh+JkPvRvvW96d1JtPj279at4KYtHgs3wt0R9gM
7UdfQuxYluPto/0dMWXIGTFqWU42X6Tr00Nr1N4rT0tjnVOObw78+vetQZVDYA+AJmueenF4On3R
Ji0KZ1OS3+UPkgctIhwwJbrBYkE1n/gOxKIKSSVtGMtZQwJ75JfG5BEK0xBiwUX8rWSHiCgY7QYI
aSk9/4Schb8rtlVuohtnWO0hznR17Yax9B2P713XsIkvrDnx1JQbccqVu+lKxidE0g95h2CSMm/1
MlUWAxNdIJSj42uQFk7QpaMuhIYJyMKqHJl1M7Y4bkj9D6nzuhDJ5E7xvUOkpt/4TbdjsvZsDOiG
7m0QGnyx0IwKErngX7uWTJ3WU8pUkfVpBIolfdysT7TYn4uy/e4QdLx0zf1CZznYNbxZNpJNUSB3
F9UX1WDu4IXtwH7/JUwMsRaqSOfxSekvhHZ59I74s2ort23Y77MSX+jiE6mQ7Vo9+yFIyh+s+dbz
a/9ueDq7g0V6+6MCgjHdZ4qU3nGC/Qs6bcPVSw86+DrZ4aOG7QofluTWMy8N1ZFgtYhESvBqYrDM
HmgTyP82jBzbHkO+/GxxboXKvDU6XaYncirF2qXy+42bxn3grq4U1+qCBVYjGrTAEkvh0MjQXwYq
4vF+K+97BFtE7rQoggAfiTmvJPQ4wP6lun3WfdP9G+dCQETJifVEOaCrZzzdnvXl03xM2a0++WwP
IRYauNz5C+p55/+AtELlq1EB5grg70dQdxsRe8Npm+3r6iRsHkafWGD3m4cDFaYgUmYIw19CUwOt
FUDpxSPsgX5IvSe7BYtCD0EtR5s1JAqdg/y+GjaqXeARvFteCuKDqronQgd9VQNCcg5kYAgnxJJt
Wygplp1qIXdoWYAdzg6c3aJj+uiCE2mfbwb1CK3nJgvmpaZqTi2HWhD0kwLCkoXTSg5FFqHYQWjN
nd7NB7GLb3T8HNtqopjHd+TWtNSrXfmYkmbwRslQXB3uHmDFeG/2mKR5WPFvdyOhnzSDaA6xI+XQ
fTUWolpV4BpPskVcR1D9IvmveRCy+cUe/0bBacKzmNPhNUxTHE6dUhl8M69hIMu2GAntdNMbXvH+
FyOZdNB1mL4VjCM2XAHgfe2SryEZei2QNPfNZsWdnLixMPUT6vY1KPV5rkUnnVj4xADOa9xvU4Xu
7aB8Qq6neR6JgcruJOanntIw7KVDwWkW2zVJIKY1IUFFlFSpIhT2e7FHlWdwNYeXt32XhU8qqkg9
WbgnH8ebbPxR3XAoQORggX4ZHYbPNpIpBC70CD4//GPqquPiA6ScHMcgyq7VcRnLI3nVHZysTXRP
H6K8l8rqiosdMUih6VjPk5pWbIVqhLSSZb1koBq7bBCdwoAAYHz3+jsL/9r2HrjjMI5ePxFWT6Pj
2Qb0PpntOLDSl1+J3E/PmizJCsqf+IsLOqQmW1L3bIbVcyhCk1fXPubwrCJpcRvuaVV+eG0C0iue
0yf7N+qcsagacdh84M5JlnKYdSAL+ptdJo9A5tXdNcCQJ/1+JeqQ/ZjgC70XGKj+oPwFReBe/aND
th2zARht6cBB6bXeZXvqdolFnxLPa15HnGIafPcSzPXUsK2GzDRdQRym4+GXFN6S4/nJ4eRfcbSX
qrzi+b03K2unxapNt5qGwnUl9KaXtj+y+sM1nWfuVO7YuQ5GmEqHy3cYjkNvfIRz04497LZurTXN
6zvmZ/nRt1aY3vTn6vzRzH8rpnl03OYKRRT8g4dsNdnrEM9+I5+N27h5AtCfc2hb4+6CfGFt+Vql
Kg12CKYEywEXsK7G/vg2nIj0XRnMxqkA042ooQRLQq6rcOesmgAWv7I/0///g7jalULsBIXXIwxp
WKUHo50C9WDLu78F9gvJQff3c0aWzgzV9OghthDigQZfiRJ++cgW400Ndv4CU+CsoEJCBVxSvhcW
McwgyE7bb3ip66fyWEBr2vorobh6Da3VqK/n5Wx7Pl3aCAVDrne/U0C2kgb5ACBYwn7Mp0Y4DZmv
H+KV1XHcELJzYqxBnS0d1s7IBl7EG4tMFLBaUsvcd8XIkp5qxT9cnXfODg7LHcCWt0OejKHhYHy2
2z7B0axq48n0qTUp/DZMFghZpvdyAxYGUf6Pxnf50Ecpfo2wO1dSHjByREqYJzpQ7EpCgE3pFmk1
r8PUOB+ZzWmEUgpiC/8V2OxQ6r6wyGJUe20h7b0CdyNHVBuxw/3gGZYyNCSPxCz2jWAxntQh3pfD
Ygw8A3HEpLQ5/3liVcPSOyvU5wrook2bITf5F/7N9E1CADAFHiUkOFh/uybFVFOR/nGfd2YO/9sb
sZS5yC0/x23fBRqqCF0S9mWSsgkjuuq6QS1JS0JTE2Gbn3nz70MzebFlIDYvGD3cUn+aVKuPRIzn
5fmx/O6NF3jsuO1zj3wgw5VevYWmerpUt797dcCPoek/r2iOY5mx3Pxgk8uGnn8pCn3ebG2rpSw9
v7KaeMAy1jPVmn4M9hgbE1pR8BK1sErCZB+0TUomGlgyaqZLLA7VraSulJ/e5xJKRXp9VZe4Z5FR
UDNA4dNzz9hVCAZXfGhucohIKxdQOkDvtvN5vCDaDYBzsRClDHXyvMkHUwUA7c+cbQv5ePT/bRfG
Cwlhd8Zs9sGoqskjMXX6KOOmh0bt2yyIsd6wnkCaiAvKKbduBgJwJdmUnnq4L9edrcPGWRZD08zQ
xgEYNnJn5CA4fVZqaWjC6qnmEVK49aaYbsiP4daaE7nNRmKBjo9vIgR5viPp5bRScwfp9XIFhbW3
cVirPqrmIIcrqxCtQkAC7DNSAsgOi6rXEToBRY8eJ2aUPR4fL/Ec8Bq93CqJrpYXFQosNqNnqfkR
Hs+IZL01nfmHMYuLO4vA9m1GLlL6O4QHFzAd9iWYgf+nzbFIn52X0JLNJRde7qy7U5nA1uZKYyVt
daR5BaWXf7sy9RRZK39YME1A6jA/JRW354rcTgGmcsTPb5NksRres0jL5gqTerEnCnEIG212uqF/
Mzgibbf42U69Est4bRDUQ0fEo2WN62NLzolA+lgAK8bluuEe7vlqMIpz6In6xRlHR38a84PPWXCs
H1WqvU9oIGQshPOqskBm53dq+IEDYebD4X7ljmdy4j1JFfshOG3Q3aNMwiFecF3go6NFREl+SHHd
0cMw4P2fsbcXdR0PkglpdlBMZSEtU5FvyeAFrDpjW+vGqkz1tGovs9F/1GrEiPHogp3Dg2EAEAd6
VoDVsX5arGZANWT76BZVfyAjuQmmoSFk9ckA0PXzM83KFO14xBZ06poHtXiZ+KxsW6tEdJkSGbIs
Owlk3NR5syy/htzZmnPEFJCIuZ9KSc3xKI7KWIXeC+Boy4dCiHkcEokIbwwFdcltZH8OWDkNE/xu
aGpBD0TQlxwAmPlgwfqWi9sRJXzF7xI4l7/8uk2mXBR+yvm+1oGQvri0wvlRwO0u0VqKi7hRM5Kq
j5XIzLs/nBWNSde+/qj651JDAIYzrepS+khkHK8+i3v5u1A4Q0ar2wiIjZsqyMdKvfwTp2mFpw+C
nSfTjFQRNb6djhMnombH/emlkLjrkpLBoyStOJenbm1DoYwxJJgUCUUyA4mxt6RllBH6Y0C2mHsQ
xqzGsv+jtdYpQL7RGmTdovFHULarVxHXyZi35+KSx4Mxgokre5lsHO+xQJBHBOzD7aoH7tU5Twz9
+2ycjGOZURoAnRZjgfavG7C2Ofa79/nbx5/P2qd+B5ifgpIblYiJfAV/FszB0s6rGMDYwMhw448Q
fjvK0UJrwujG58kdJPmgnMHUpqw9TvuLOaQvn6GzF5Iup+amrdFCASv/HfAp3ZUppBu8zutkhZ6s
C+fGMAtU+s29Luf4CWa9IFwdey3xAjnr1L3kNDNUIEHo6/bLFBTn2B0Y9LtmH1iUregmZy0Z+s19
egNWhQfokfeVaG6Wt1gpgHXP2OKxF12TRw8HCRP2EgW9D41pY8srTiyjH1bgOcGEZCEB3qNzwDXW
tZHeON53kKbEolek9wK0gKhWBJiPccoC5YDxguom74jAVPKFpYK0Bx/3npfWWoetjK3ZNRVSZklr
3UPgWYxcY9VJe4bmYJyLQPTiKs/fW/pHN+phcDvFePX6fyPqM2EtsmqW+yir8xVN9fSzH07S74P1
rbZCzOpPv4o2bjdjecl81qbDHKfSxA7muWJmhqtLAxGEUVVe8lX1VlPiD+MBx1hEQvLwMNbMS5x7
OvO1rNmoOGaZw9/MNhaSfqcr6WvlMaNr2LLuFP1KbrzmWJVrhVJ8gn/0reT0DSEAaoD5wBcZ/T5E
cIFHd7G6bUUx1kJU0+PTiH7qBwz5QbvOReFC2QRn/iJjFBzP8R6Aga+AmHPSnQ34iGJz3RgaC2W4
sUV75dBd8xFwDKwbrN/QVupk0neImEAKIvBhrP312sGFexjppYBQv8FnYjYr8ngZg18hbxR8vr1U
RM0kGxhPZrLnOZKtm/8eD7z42qXmoOyQUVhLDbMSA5XNfiAl5HvMv+0CawcBTxN2XM+RRSG3E5Ol
jLCYOUgd1T6Wl4eqXWtFH9hqVyA5gBqQ6ScjR4KruM84RHY6Vc+gQfHEVZXILq3mX7quQ99W82Ce
lWpLMqdLrHD3FvXOJlbFLL3ap0vp0sMkRK05MGvJFlfv+5Q8bFRjFJU9PPNP4tZckiDFZ3Tgr1bd
Nio3HeboQkQt+6XIeDlHYtX+DjHAETwMOvbBKnqWAH7XAAB1MiZ0M263TLKlTICkviLYexQFM8Sb
lpBYBDU3Ah/AkCk00hJB6JTnP443gVLQf/lOatdiAo9+bcSMD42KBEU3difF0ZAU01wmhFjy3zSJ
donA1swD7jixfAT0dS4REQ7KFZv5mwuCQjK88vLol4oJPN1Xhe2GjvIdxrUlI9XMvLoS/f+mrFn+
+1ichaPFmPrDkl/H+ekqYyIVIXQ4UfpztQA+akF6A8HGmxH4gou3MSRwbwMZhSt080srs1iHHubT
qCYIsj79VH2UR26Or0C4HZZTLXuJ6Y+8IAs+4bVpmwf44yhYPdiKMtIcnMK2fIIt5SckGqez5RE3
ZBTAAwkU01cRenur/KRjEWU0Ukq721FwXL7qA66q2OhQIW1B2pBV3DBIMTs5+PS48m/ClIXmQSLY
UEoHL+2eNe0AqlRw7xdLM9Qq1hVIiM7AHY4vbvwWxUrylNYWAiq1NXd5EiHWPeml8MfiRTSbJRTY
XNs6lI+ttDeLZ3htliYLlR0quNiGSrujEbC2Y5+tsj9iKRq5YAn20G6gAObwAAMVNroRlxaCkpFk
i/n27fDOKu0khZfuzWp8j848oyOzrcAx7GiyHe62MfsV04M7VsryTUSPU+C6/i1jWhWymk2EAdPM
PUlPA33ZyfNO80DC8Xld1z4n+bFxM5yE6YsYPGxoMfpWXCvKCbKN464/9Zz1OkLkwngvCOedQXqh
xoS2OHBJAbknIerqDtEdaVxaOs111ftIuWLTWM5CeTeL/jFQ0lKwfeyjLOYo/bhh/BXpCK7JkFOB
jTbmIFhcRfIkuh3+FUfm+/+aWGYktbInBdr2PxUbh+Ido0gWHpBsyYKt3hnvGrtAzEWSxhipFz96
nkb/7+lVN6Q1L6VfuXi5pHXq+hA1MJPaRBrjUq2kbWCg/gZF1Sk5pVI8A+eb9qmV9Oqm+faNpI3l
SVYD1JaWabkumH1NSlNIz1FkIu1hqZTfeekcPC3Wf0n8OI7XAwDb8ztmEoqDjexg31QmjkIqgZ5P
tKOWLh61i5mHJyRi1XAeIyKpyAwPNc/emaJCfuzSHK5owjf1MeGdOLKS1fMwv03Zb/ODoF00bDil
B3HixCmciLQDfMWpmYtM4ZwHhsyOHGaNpOiDawhWFAfpLCWvV3UcwANbqw46jePce/sg1ROTui8i
4EY7Ug6qW494iOhpfsVVQnBnDvahaCIIcqKE+aCZJEHGGHYOLe6bEHg5g6l6pp95P2297PgKhJfS
wP/WrckI1sfhTOob2PUcG2BCyo0tf1D3MjZr4gBtFFe6LXsOnSPOtbh4gBUt4UcDlrrfRDk/N/XP
cuQ9yo2KI7opzooxPdaBcYhLgj2WtpoSl7GYUArWQHDdXr2mPV2ukb29F05EMUK3jkbn5WuSzHcX
yRiZGHXEjMJ6Zorsc4dEGwQTyUU97P3PUIOq9WkFTEEbeoB1AWkyuJMi9vadbOlZDSef4+KBw3uj
8lsEtCLl7wg13mqK7A60J2u1IG5fMRM/6uJMrb38929zPrSrD9NoaWOZkuJ7ikdqf2sLhB7e2k7Q
gUbT8xN50dZp8dCYiOuC9xm2GJBLWKVQSdc5aJpbojYo4bXs3A2gf6/Tq0CcgNqWHHZZGo8bNqET
foDG0VVuDy/IHX5LXuHwKTMI63/9x3BfCyNyeMgzAkNDTrDMTF+q/RmkTJCuK/RRI41vinUzrf0n
sy0/pETJOWoFjgnifDyfFKmeMJP7LPqkFFnurWaDrJj584zvYV7fgLiEXMy3WtELXpTpX2J1tPtj
3cp6q2O8j4rsHRufHimIZvzS433JyYnbpAqmlwFdqK0U1w5W75q84/xn6yJMuFExlBN7lRd/iQ4C
D1gmiAVNLmFP793bTkVPvr3qu2FFVRrWGFHj2k0ySQ0+xGdVybwaHPweUsNheXGBEuIGuMHEWTyX
a6F3lFFfAx6FgHaTw3XYUR5VsdeAB7Unrg+WZNSCeySN0kvaN9hbok0ChbnwselPSRosiNqcmljW
km0wcpwEoTSXFuHEcFcyB/wstz5/EFB30koi66yXwAcxseGcgOsZadn7Kt9soYOgo7H5/pk1l1PB
ReydyA2eS7pc+lze82nUH/eTmIG5S+NgPUQLxFUme/aWbQ9yLyA1WYLD+z58TpligLqUjxhYARpJ
ngNhwTsmagN0Gy9wjKSZiFzJqV4DGN1zGeABXukLc/MUcc4GE6iECQqrTucjhv6bAIYoSi2/J84m
/VWZ5TIpvpIobBNhSh01npz2bPLqpklc9LRoqZzRDhxfXqA7ovMmgGj7VdsfBm9TFOsLzouJFDBO
gwGRx/vyfpINVLQGszuTP0Ecj3Q1Xk1Zpv/8PP5WTvk+S5tJcZkKdPpUPDxVF+z7PAegTicKTTDQ
ASGSzbd6zEVC69e5V/ciFD8XmTW9o+R4fdz2vprU1kA3qcJ3/kKLccjYzGWyKIDYPZMzAmJ0BEEy
l3RHxcMv2BHq0hNl8bNFK7mxtOpOSRdEXlX6qkXIoGe1kCsz+AqHPguXaifWdHAPDfNXNT3zYqE8
ZwEn2tYDmceUVs9DlQFfPSEmeMlS4eVk2eOzcn+c6xHhfaKZGX2U/ri5wx3WnJvb9dPkiI69VZEn
Mgcb5N/cdF0IM/Ef89ExEksRLkJ0eqQnZ7CCPVWEL/0bUBk+nVwZYFh4K90+N/f0On0DAM/3oEsr
+0UQqb4RgS822O62ujQOgc0i8+Y3dR/cn3ED9yiBz0FSwf8HrLZuwV82z2fmZXsDs6ijfoSY2ROK
zzfKaX7H00jzOLKsY5+7Mb+vOZ1EaFDYa5LLap3GLFQxLkOn5YTIiGYw4ectZsxTt3XVExi9aMkF
X+3mxIbDXQHMBbIbAC+WI4goe0ZzxfUmXCuu54DSB3AEWFSkvUocyZY/qdmH2ouGXPcfSDpKpr7f
Zc1M/2BCEUqezU8ZgKtIDi/us+f+vdTVQf9m+N8LaLv02kNfGuqULaaNWsgc5z6mvzPUPU6dfMWN
j3uB++d4Ma8b889ZCU3n1HNulB/5YH2H79RkMfVsjRHQomLaOti0+mkOzmWVFx5mUz3q/FsAcyfj
/tuyT7QY/b+Xrae8AiIssghcmGJcolk7MljmQOAH/FVBOAMMT6j1rmQwCggekqVRmpN2FNAF60bp
9FE5bnyEkSIJjugLiDi7CprM7zToEN6PwDTsR/dHhPtm6mWZJD4EbT0geDQ7O3BtrisuGY3EAeGs
DQzLuGRZeMWTLPWQDwSaaqJyVRbypHANA3mSVQYihNZ0gu11DwJP5n8aNkQRcfS9y2YMhnnfl4pt
/p9gMW8NI1P4km3k7dVVjNK1OrnXXJ6OB00BjlE3dMzsID8oPwZQuuGxsTLtEzTu4KzKLqKzB3+G
WC6z32eSyNgIScL2jnpqHnp2dtcRI+gX5HG9cUsO7Dtv8syVmTve8w5aFsq21W26f27eMl2Mfs+e
FBRszM+7zsGw235VjioM/WJk9CXK4HlXDLqTgeIV1P2NGN/kx3QP43X+Kf8t7OMe2lnDCuNEXnSH
KfjF4JnuUqbeGwTrEymKHYFN7KFXBZBIMI+g5Y2jt+9EZ4FuEj1dzu0HgwbKv7rTRVrGLvDdWdw5
lCA/Ggr/YfI0em5JUBQF+L7siihRojNVHLdhYwjKB3mMSPWwL+dUVPlivEffulRbJ++Qry5oP1yc
naZj/N7Ds1yUWzfI4RiHoQLKEVJnH9gxgSkUD17jMxKe06N4VbNwI7o64hqPGeap566HZKfE0z1T
YqBfXNphUl9YntpW7ANjiH9xTlpkdNPA7smmJtek1/xy8CclKJzBjMELNlel/B7PV6Yq+YWfmsjY
CDc8SXQpMTILFFG8phbNXZqyPyQURuMn2StDKb8ZfJoiWGM4d3J5IVJo6VZsUBJX1Rs4SsLMAMXy
AK2QtensGR3U4JymN/K03bjlvzKZysAGRshurm21psgURl1Z2xRY+LAhspSwWvwyFx/Yg+tyePK3
b1wA6aP8yiQKoQa6lWTf+bre7P+GGWk6CD/c4nocHHYuevxGVcQjCbMy0J5GFOJ3S2efO5euLA7R
YTEs1ajRcNLycjS0tzDiSTMdHi7EOFkrAgdrk8F7fdshZtjig73mlgoc72E2ItibbXvbXVPVo1mO
DteoeyAI5SVPjYayuj1UcDP6YYG/t8XWbgpdAZwLQ4Ss7FxMD4csFHVh6vzI7ZF9Aw0aAuXG90r0
TaEUpoA9c/6lXiFWOBcF+bXFEamyjVxGz1kc6fi4heJ7HV2gwoayVWbA9sSoqTELCM4ew5D7TT1s
QiNnPA57vRdbbR6br7XEia5laa82o+RdvH3JUJi7bSf/Ur+6g16vq5JVyF3MUi+dJux/BI+m++aQ
JDPyHn8Sm0oKdX4ZBZWDpBTbBdpDNZmD+a3H7I0xlE+67whn1IM0WcYW/Tc7UHD2nBT/56MPS1Rt
x7kvK1tefq8vdkFSQtMFWjyIMwdGb0bCfZLSDMRo7o4/WGnJqOzJ5BGFaGC2VjDs0/HNBIjaz6o+
6zLsG8043Pty1IIUfrxZa330KFgNA6Z1qAXTSKZZfkmx2d7mLNkd/mER5/JPMNxT4lX9HYvZh/ZF
y1xyyyPsCySDqdprmm9O2dlZJHZuNw85NjZHEq6tFNA9GnoCrA/5R5Ad6rFSVD9F5ILlVbAqy0Jg
YgmkR5DSf904dc5QDEx34rbXjtT92EYG46bjpuIcFtkIj5AH4yvj9f//hbfBOfIp7qbvH6+OauXM
elbfFbta6s611WxLFWIuP8zc5jbYtl231Lo6jYer2zJJALG6OLJxSNgFwZJfOe2KbovGNBNux5bT
XwnmQ74f0cIGalAb2Eoc6j3t+tD83rHvM1SMK82KBOqJFBVgzSptfLJG5Ky8ECi4tDZXprh3Es34
INUQDMq3ha9R/afL5YtlS3UhQS+zBsqE0QomHZN2UVGiPtyQ2tJqklJo1S5eguiEsHaPqCMIZwxh
8romFXUKjq+7qQVbCg1xtSXtu4ND/c1o1HIBXxd045rwaBjU1uDAentQwuQAQzaYWcuoYtweIAH7
NPdg4dEHsT9SMncXFIvo4mMVNHOypTEL/C2481TAHbbgjoC/epmJ74OLqKEhF0uXhDxDdPvNwG5U
ED8AGpEzVfUL6qn7bssJhPmDIcqHrQmZtBBxnLVR+RMacwpv+JgMCgik9eyFW2IhjP8T4qmcjtAj
9VIblRD4lbXc/ArER8Cs3cTdJXPbR638JxoVdjUTAcUSh3Q58MixxHPB03JfY/3CxCR/jOvwLozJ
cYMBaahTQA4DOxyvH3GAPyB/5JuX2aw7AfjSDRz/aTmtzfBygAm4DrU2V4dgriMfXkICJyazde3m
McEWad/dyCpbk+7zW8LjEtg3uQlfhsqkZF0bnYi36/OqFh4jq3gO53MKh+qqqjdiEm2ApfTpw4yI
a5qSME2SozBYUbHkXe0AMAbzAlpSpNiQ7ZMM4zecVMQyi2Su+jE0Z/9vhyLbyN0etzO9md3ydBJA
dnIstBdE5rOfxPej8Zq3NJ5Df98vP5BHqrj2h7E9tzeaodzSoSztuxurVVsZ3LbSz+3NBoRMloto
jhD8tz6Wdzmiln6D2wOKqg8kHaoXwEVPKmVIwFWaWgl9PoK5wZdG62PD3/sQ7K8pwkqQR3Ip9z/6
4HiMj+tMyWs2sOOM8FXPdXpYRIY9T/P870CeAy185xm4mzLwVXhX3GwJvtlz2pSho7ekBNPkKZks
a8dQNSjt9kpReVpy8tVxxX7UYaWrtomoTGczEP5daDy9tfHsnk85VzCfs8bZYEesuc1emZQUp1HS
aXPDeBVicX+ZJNldKj4Hg7NDl4BkUAngrtAdouY1vGrVsdCU4kus3ft9S5lGTmJS2O9H3TiRkO46
zY2QsGM91naWixTQlA36zP9/IJKKxdOCBAZTnSmHhXMLJmoNTGT05qR5LZVG5W0Y2UzgJiNO/w1x
bt79cnuYCKyPKeP4pSZKijHVVtyxdLbYHG25wNV1/cs0wbiodJkUme6k6WJ4ItA+X6eTkLKUokP2
Jo9Gudb/LJx7hW6FClhAFGIns1iOWeNEJxaDvxKA3v+z90fh98109xFE+8dWjYMo6mAIGMG5bAhv
w5SMF26HRSmX8rTk0i/3APqol4u+nkKcfXde5ZWjEfQD8F19tT13yKaUbhKu+xA0JuhSSJFOQ2Qn
LS+RM09C3HHSElXUg1yMLZFnH0XrBmCCSFLQtc2EpGu+0gL8JRUWPefdDarODcgdydstfO9cNAj+
Pll/WqM1D+LPFSR7LkFCm28EbTARswZLWydTMeK7Oh8fmnbfyo97oGTB5COtyCT1hBNryyt4TKZC
yEd6Xp6Wm7pQz+8IFG+4cZ580Y1uNBPiiJSbrKuZB/+NSHN9JVyW9lVyIVua7pNSH1K88Y6XIS4z
b+zmJkKVwISUCbswM9Bez33h5vHE4QfF+dOdae6M69QrGaHBroQec3SJg+7c1dSo7POHpMIlbUUa
gIxlh/ePRJ6gg8OyEjjgdhnySw6uvQwQnoEhqGyMOczLZmb0olHf1OqOAK1IVfR5p1wZpdVUEanQ
8iBIw3bBCWZv3XcA3sVLh5pQG/vhAJa41Tm1z79PJ3drCqyY9kqy0pv5YACp9zGr9hbcHJSFVA+T
oxjJ38rKoJ6eJ+wi8teteYxqd8R5Odp6MHb5SjhmHT4ce8fMxGccZruqax4zBNLpMpsBrRyn8rNx
pAkolnOGSC66u3TGtKZegtbyhrASspj/RW4LClUPsazZgpuPKp6SQhw0XyuIpSfdsXnkgH3gmmKG
vf0lnAaxbo5AvpmVUWNlEaLE2284IxmgF2fqOSVnWNtsGF1CihaUhj9RBycDVJScCr1ihd7UjB5D
mMA4VP87VNtTpaEA9V5Bsfx+5mVEXRIV77YzNSlABfG/qeaFKntcQtuc5Mx3K6ORUMZOboio6LoY
jPiJxJ8QLmJpKIZkO7RSg35Mq03pSOuIsSeMoVKZgruB2fOm9ymiZ76VGr5NCQZLyUJMQ3Pwco2M
PA2cR4c4eABmfVF/mIiJTOcy6AfKXh/eUjSeTQO0w0V2zQVx2wD2L7qKnWuqs2GF0MWL5kFcbrhA
i0ODxL3EjWSTtSLM3oA9/hhjFWdCQZtHeRPhNLa7jL8jlktJtoF2Esxmp1bydoZOHD85p8q9N5Hl
VEB4PYdUElxfL28188eoEd806PpRV/jj1S06eA+u3RkZQs0w1209f2rcqf24M2ZlytoVtsl1gpTN
LMR2xWSmvDrTW438oP1FJyC3NHKit7ON3efK2ZVQZrMaJ+LqGDZabRJt8s+sZOCSNZYuQvm50ndw
kq33RoPEvxom0B+s354Le4UqZi3w9n2Gm/VVC2XPqt8WMlPHUk7XpALm2MMyOLtzOmw60KVPsg7/
TlkcRuQizqT0QKuqluskFzUpBNNWccWf2A6DD6rBcv04+ZAHgcKuqzCk7mDfD2L0bH1tbDCHVOoI
CDMyt+DMIEnDmDLHXAGA5+3mo7TIJgiOroBVuRlRSrjXj09YBb4EqOuItwEnqoSJ7oV2oyZkJzct
LUM9Xb+gg96utwyK5TJwfsBa1AGpktnvQgsFhQ/tXlyEO4lLNAzA/ZZE9zIhNPPhZm3rBQHdTKcC
ot1tBMVdW5IKqFrhGlKecjWHYkoTn3mIhXXylKqFQDXyfQ3L7uyEfEUQMU+9zc/TBZwO/GpBBHre
ycjal+0vsziG+tdnzjjqdeWJ8EQOZrk539aY0DgjrZVB52rd/5B4Vxtuq5kiQJzqoqNPLEP7Ovsb
85EH0UEpeaNXxzLaZULeQFqAf4A7EICDc/Oih/uzgDZ/D2M4zDml8xZAoIz+G+H1+f29U0L84mIw
dc+13Xzc7k1iVCY11OX8wCbYdkzr9KJdN7SkaS0CD9b5xKiUSG9RdKXcfTu4mO5luu7om1FL6iqI
2ycHJiWZExH7VegIn6zp1Sd7L9UzGCIakwF1aR6/iCAmqStR0sVuFKTBzYKsZlKvaOY2Zadql+pg
DGomMWj9mR0/7Tx7EhjD2NuR7v4Rtmk4Z4woRLuuhafsHXO0JZ95nZOZdF0JrElFuVSZQQbIS1mJ
J05oRMXTIwLdfPE/bYVPnJNonbtP/NWgo+Sb5rL7vKY19zsXkc2pk6J+EulE3qpIsOkb0bZLeyjp
AUx8RriJLgReCL4aGm/RfLVk/QUK2LjDdyjJZmOB/750JiPckvghFWydIgkB/yvq2LSaT/gZohv9
3AjvQY6gKzkTM1/S4LBE3SO3xHCSk2lq1XGFeJEb/BqRFPDQEP7GZDIytfrrJxbYsEduz7uv5eCr
/v0012gj++ehnblCjoenPo6HrD+z6/eyIcH6ibxhEqwH7GQ7vSf4B/z7UvjHiBMVjc761UYJlMlD
V01e9+uENTHQ/3raVbuWCuUHGdpVYnzggeIqNoGtAJOWciaB2+t24Gg9gw/OFclOv61Od6JN056E
Ngk2fMyNWbnLU90lX0K7pccKHTMEO8fvj877WymEIXNzdZf2jLFlW0BNFFKPr1dFQxKKvrVCoBiJ
09HkgCVwIEsLiNVvZNUmMncTC5bbooxMTl3+3LSJ9YSZDt9zLT5doiIoK9nUJMi1ZvAQDe62R5GC
A7IS8Fwtu8n9V/X2sF9UQC5mT2qsAnPL+4rcxfryjvBl763LJeHumqcmbeCGHSU7EwGXfZckVgKz
Tr71umFfW62g4ZiLbi8Ou1plG/Qr6oxbqR1F7QlJgauJIZyWyrezRev4L8O0Quyjpu6uCQKImpMr
5s3H4KEvLXhXVmgXu+03jkW6ytWHlPS+NCm7ByWsQUw4z+ArPt1uwLODDptlQOktrIeINPs4xvRI
8nLNjqj2IevS3cUrcfL2TPxX5iJZcOl764imhmGd677iwC91gyBfFKS7BQeEnONG9X2gDxd79jZQ
NDSPwH8uTkM8/9wNxCxyw5BQU0WtPUSibgczJbRxQiG3c03+NrGzBYt9ioV1lfCtjDHbOBbd8dtS
psPebpKwIpg9QwuZas9ibSTpPPEJYkz725EIpTqpofEOgyOC4OlqyBtv80X4DGhvic3ibQjjY4XC
EZzhBNrKXdDYNiIyIAYbNcuDhk68Byf0L/iWUx6FGZ/QeQOYBru8u4KYcMollqnieLo4sZJjmxsv
j/GajOPVgSeQuNbM+1SXWyAiLLfTYTx3fh2aRby7lnrmzOJ/pBhBdNZ/sE0Xorg2wRC6kUV3MRyr
1kkkIfiPPprncKcCHEbnl6/bWigPkapZXQNCg4L47bPb3qiVp/tFjXMteCGUnEiYQWCHqptztXpT
idD1BSauimXRKHD9Uhjrg+fPR8g41NxCkZRWwu2WGcKZ4t1PRxN770JAgZASEENHTRdQeA7AcMgO
VsHxZRiShC3zmOd3vBWtCmNb1Jlj76znoegIKzvfLpQslJrETck9zis7BP3oQc84HFa72vKW6LEC
/2wVrvAw31dcmmbtOD0TkYwoK12SvDFVYexzgBMW/oAppHMq+6cbLdL17OtmXx75CY+NblpbdvGv
X7bpRhHdC2D7Gc74eljrOZ7pGa+HSj7a+qP3HGqV1ueUFDN5AZfmCyw741ecLLxVmcVI5GzIoMKn
xVVkoHnBZLZ12RZzOqZxV/+hzx12jqiVIPTrfq+zMP6J/YJh3NyymkIfegduGpyiwGuOt8L1UPUg
X77rURgyX2O+QLeF+OZbFO9Mk2L2ZQxFokWzAuyOsv8712EDS/ao+Naa+jDH0HjNTxyrEoZHVoaO
+VFeTUeGMaN8OfIaX5Pr1Vk0LhwZfWOlL+/eixbGxPNGv9B53gtdmKlTzL+KZzrwRDgVDlPKaWNh
0hajxZtCfUjGn4NQ+nQd5EVwnYdIjjvnyPGeYmgF9HlzxZvQsSncQDJiCfuFumzQcDuBWGaVoOJC
EzxX4u4bE5lRG/gT3d4IHa3bO9nEkhVaRHvMY5ZuowejM7NPzhELb/L/JPxQAAbLfNzPbOSQV5aP
SqyHaRj5W4HYwL4uF5VO4TJ/p6ctq+DUJzFwyXF2Qa6zz48kXGbbcHak8YRoQWLSCSaIztgYJjlv
C3f0gUZRmrT2E8WXp3UpyX1dDP13q3+EsINFkb61wToKoeeM8jFjC5GvVTlkTTS6BaNqeVrke4oJ
bic/mNVnzL1Tp3oZDaPUpE+TSLQ/F+lcbX+v696Di3lx38BwP4Rhj3uRU9FatMtK/WXfbj5IBh6m
iO87Zf5g7BqOM0KA/gA7w2rOO7n3eMMrqlNnSp25jKtWrWxMVbz4XcpTrVDstmMlaV5qJOS9sy3C
ofy/F8vce4n7EayBelmDBJ/urpbM8W5jSmTtjKc4isnQKo5yODwRi1VU+IOf3eAOch8ED4suaM4Q
WxTSL+otkqgFoVBi5q4PYZYtwtcfeMDettw266qhDE5MK9yWT1k1y+mGx9XD2FTUucYbLQf0+p2m
/fimEGLLGZ65yalgjE4Tarip/dj3+PflDzFBGH/7q9cb+L5B0ty5U2XoWZPA4yJ0sZG00O69Ldyu
0VDhxU7uSG3UqrMqYIQ5fpCm0oqE4AJjoVlbLt64VSPX7I9qsB7vNZwq88kCAgQOD5HtmPR56O0Y
nYidQwKzPpXt+YGXXbofp+H1pGuWM8hfvTmmB27dvysCvbkVdXXGdLrtzF6GtnC6DHQ/clqHTr9z
W1O3okD3e6Lys6NWGZB/HrhT+PCkD4uybILD9nOAu9i+FtjzPhdxCXMM5v7qYSCtd9209zHpOqZg
r+gryZs4zd3DmknVLPIuh1QDxc9tqFKJytCa5aD1aHtnGsX2UlzraNPoMVx1X1djRzDcczY4eV4K
6wXZ0tb03+MGZNEubqdbM1jPBQNtSgWfL3UTXMoQIK3sS5yZMpbHnPfh1ef3LOpt9t345L+r4Jjp
OJOGz+EkRA7LGa2BGK50/XbFblNB+4gCeIBE+Q9Cvot0E2oTeYsnWwOtZr0k9Wkoz8APn40ce/Xe
7DhFIQIs6mc5VZj9thgoUYgxmWziitVI5mxXoEc+sLyx/abqQJBjNG2NQe3PoAgIGt8BaxHcLwPb
UeElgumGh6NFpJoKNpz5tffYxQCLYNnuOepRjB1iuZvj93tsseudBzNOl3ISAavHNAhoiJOM28+0
u4IMXTVx50gM1E4v8RAkJC6ecK0mKHBvsp0wXIhhw9jWuSZQs/898ConLy+98BeMkCl63ZOO0hrg
GOwOadbxoF6K4rF4Ckncc4bQ74Mwl0vkrL5+aaOp/DRMGXwxhYGQngW0FnRRF5Hu1sXYgOG2vkkS
GDqb3lCIYwRWcm33zZSDixXYWRw6TpEBJBkgUtjoSk3DQ/RNkOfENucsQO7ApKjypSlC8RUcJ7PR
/wXHo0BLV+6FVaVDaX/EFCIeKJ8PVE1j0IoPJJ0cJZQ8Klsy7OdQFOLllmBfFVoHxAgyEzaD1+VP
qCIHWHqJTVlQD8fzzibcYOf7xfwG9oXQ2q3iqdT/qDlCpK5tBUk0CKvZ0G3bzgViSz/ACgKGDTSi
+3xbmgN+hJ++wONcLfeiphMCaxs2r0+5RUdVMBoFMmqminavx4AN5sK4HHXN/K3vykAr1UE+coGX
B1SCss0/kcpSvanxsRS9NX/f/DYEiQ5VK7397KY8DrQD1NSrl5VYbGrsbGMX96Lt6SCEswqpa5bX
CNMyT2S3hiq0MnWBNYD/JTyXClrxVnnZpz6Hhhc90N14O6NXBBcTf7dvRJnimPgzqWEJpjCrEksM
3I4JoDZel4Vd/+j1t2xRD8ii19rpylURKTb6na0HJXxAny0vDwyhEVGIHf7tkT3HS8q598S4s3Wi
Y5CVVvWqcM0tv5PwiPh4GgSEwKWn3VR9kGWdE4b7AQLACb7lQv+4dN7fj/89fcvDLnJcNxKlAkPt
YhwHLhxAhFgDD4uWpXUU/4nDgljCbIi3jnXnAqqTtSg6RaMaSiHO60pDb4ot2xP9M0atwBLmE3m7
9zZZWI2e1IbatimKgxhaV2+YGi8++s/RROAAdjSnzy5E5CCvwSpLjMTSagKWBav6Y4EccMo08i9D
Twl0/xusCNZ4nsvGpUDxUI/kQiLPHl4mrGeOOLRCgT4gil8L6aLgQ/VzjZvJl2dsqC91cihMp+0D
9Awcodcsvkn4mn5blNUr1wcf8h4dgp8TM3KU3XP6FSTcN2u/ifHpJzFATbgGqc1GcnlbljNU4vnT
M+fWtvf4jm70k0cs3WW67ZHrfpNmDJ96PHsYQaXihtuy/ZQ/XMa2lgP9kPtmADEUA7pttekUn3Ma
7Q7swxUA5N2N48nJVWHmCUoKU/3ap5nO2vHmWbJiYxfFdHGdj98zCu7ACIzI5nPNsd+9lEvkADoQ
/cWLs0swxr1pCE7Jp30CUHNfAJgh+x7VE6PQy0aF2IBebNHf2LThFuZriCDl1HIJ95u1AdF0XC6l
Dah7IKi9eQVs5wcB19KDle3hykVDPsKXy9L6wZQNkK9tUL70wNcm4U2fMgXYOLmf1ywRjDYdBK0G
t03x2hd+VZUlKO1kRBZQjWRrOaOot7fIj6e2FXXr00/UDAzzAfOWR2YFDom+ElKsfHU4MY/WRKPB
hVUsK1VOWVXoISNRqRVSUw39cc8qtPwcaq9HtJpMrWiZxyRZiPgUh/k2EsDTJznO5Tb4qQlPf9ey
GrWgyu9TjmBPLs8txx3Blkn/kLuG6h9zgHNXSwCOg8QequVaOrDX+sr/n97/JuRSq21Agg2euCrf
nxmnG0iKkDf7twa/7MPST3kPNivaMcx+Yzp/oGJeYxW4Fpz2BpEU+E1t7iHnqybvaJyz1fiE0Y14
vvqqsu/LwnVmIcfQUOBirujW0mI4vs0aIf080sf8JY61uOCM8taqf3/uKzF+RX1QsvSdMa5TahHZ
nVO7TPz0dqR9a/O5RIICSWUizjRtiPNlf3OldpnF6jeKKUA1If7tgmhrkdq8fOJp2NOmy9x0re1x
LmOZ9itAz+/VtDZV1Zj2JE51czE+rAQxNrPlF2JUTWbPMVtBGPOhpMSjU2VwtfVEJ+y3sKXyeyzT
co12ur0x8he6a2uHYc2vZnyjq6ubTkrWT846kdTmlPIspXDY7Si5p9v8jKUThzqSGWzrM2+7ugqR
wpoiDbk9bGoEa3VfozhVphXW6mqxpnbSOGZKbPCsFLqbw/886WIRmQx+cG3YAlrgB4MPR44N94aY
sqd0pcMdZrp9VHdu1Uc2p+JfWwD1p8cbJYEIwlxoJMO4qKQqw3QIVWN7ECh3Y+6F7/TL1y/usaCS
pyIU40dP3pSVFNJwVKF1cWs+/BkL66XNI5gyLgDI+i45sGghRjoHh1Xt/BV6zyMBOp6h+q559f3v
uUzYJS3k2eLgCgV0ak8YcJGs2PH5JT9/Mpc//uZQnV0OobSOqW+Hz/2tzOy+xj7lny+X+6Eut45f
V6y6jdxjxp9HPFOGyOVoIQXQwKu9Wf9txxpD5Md1aRnNb036TQj/AiLhGNeFD37OVsAGTUqcKk1H
3EHeMr9CFs0o2URWgl+3wR9/k2rlOKuItYigT4hXAfXtawTKhxW+NmMvFgk+Wg531f5/RaOlE6Zv
hddAvy0sh6ebxx+gWEnLWR1VBaFI+gy349vUxMi9ZDgSB9rPyCTckwVEMrc/kxExXqdZcZ/ghhR4
wuXS+b4QSMIrRa/EyF6qzq/9ageDo0LOHm+2mtayTRwaO0LKPjs3Pd/v24MatefrZxv+aOj81m10
XWMaevOxYO6vAayIruPGZYqcl2vIEOgkZyhWarkMD7s7NkfkRMQeDYugASfx5tOopBeRz/NqDp+s
HmD77O3j7Xlj2RG/NGotZTTJhjbaWT5w+LwnzNvaSKCuBvfytSxTU1XKkt1ki4DTWA2XDUnKSR4o
LM4W0lRIKgxIEfPYJzOqY9aTrieTPrO19sjdV7CbHlZPOEAH9uOEP9x1Qwrrz79r/faZp3IEHdlk
Y2WTqsDQ2R0RWPNCYGLbsAJ5Z/ol34EaTHqth3Pjr118dhHyZgj3Zut3qXKhtHPodynZp5Q34wP0
p3IibyDPAj045TzBUjSnovekLEnV34KPhMbUUY0bjwOuK813L0UE834RDCFaAfO38g01zHxQFGkl
0C4MTY6VARm1XdvpW6Wu9y+3uQ/7n4z9kTNQ0EbYG9v2w++GbQI1PfOSI5RwhZvAWL5zT4ppPv+s
KXl8+VzoA5yXdkQOFBU9O0WJ/0qfUHDHO+x/pngZWzFDE0j9YVCTHAFi952bvt5I+FrdC7+WJRBf
XC6unzHfskiGANpQwJczpsjhng31+AT6h0RMVxuwKXOAbZ+xgnbnjXXR82d2LXlldL6p/zyH6tWE
FOBh0SaSZ9r4EZ9cgOC46wGd35i1MOO8L1JdwtMRBD/A4vNn4y/esPf8+N2AsOQEtzIFMnT8EsFq
dvoTNNhiRstB0BTdadkyz2j5E2BaoJUALwrsav4GhD9ti/LUns65zM2bbDcMQgKuSCabU433W7s1
4wdfnaWDEyeXQCllrN9ah155zENsKNRUoNvq7HLznTXez+2YcI7+Cwiuwvf70aAQYLMxIjLXEmUM
XrLS13f9QT3wW+tjztXsL0efG9m3l51R0fssandqur8ztvd2LIKmxjEJo7WTF6MWGlFDbBGBBrIS
gEfy1EOvhsiySdUEe6JHH2XC5qi+KYk5kQO50mHJrXWoJ1c7eh4Qt4nlRw6q4js04UtpMemkiEV3
9PDPJpTMKGAhzolNDiHmTbpy3Pmz+GSHtETCktIBi9dPII/uEopCkIzO3AKTs8mwZLn6w2YHiGQX
JLQ64fLBiZPFQpEBEctTowhBGzpjpubq7hzjvbCd4F5egTJfLp1/4qtwXvhcYdnaxAZqRhG/+70U
Ebh/Gx6bYk5Q68ZeYlbLFuzwVpL/r/6x2pxnAru66oVuNrlmDvLY/S4QhmSE8PvLZD6/Rwk/e8Lk
fxiToMN/Wp7DcYQXSV06nuXmXX4YQgLtfBMHCKi8lIpaQEd0H5LDnTAi4CJkeXJ1UbqORxdW7fOc
oQr+W/Zb0ffYuz7bELZVFj2qmhgWNrOFZhHJuG4IBfZ3UYL//Zd0vOTcAbAnG5Fbn1tGz9knkcjR
ozrS1HZjbeDoi+4ucBh1z6qSImCdTfafdZtL54ed3YVZEVMULJFOGJOut2xFEU+g4xaOOE5RKo3t
CO8FThH/5Y4GTaHQ3/LTbbH5LyXz1Vc1CpFXc9meCk3z0OLXSawrGpu44D8O8+Z05GNtL0VRN/Sq
RgQIv4+G1xqpi3N7XXuT3gMw2c5am6WBUuwRYMq1egEBRWhmBaVYxe4yOSBSNpei3gPoBpDYXAc/
1IcvNYMkYiuaZfj5BfZp9zhkp6Utw2bk3lZf4cMsJrZx3kqhboqP5yQX1IVZaK4baW739/Jd26un
eLs1X8KLgH9scpnRfbcc0xDZ7C3r5nsqUZR5Dr64pjfTzn2L3w5bTL4XeXK/09QyVPOg0Paq1FKW
yzo9s8YogGFV4SsFKpAn42W9StbjsznYhrq5dE28hHpG8fNWqEjel/mSlbiB11ecrOFrvhq5tCpe
BL2Jk5A1Ddg4G+oGl43AIl0wqphzKa9X9f/ci8CWgTeKRSTpG8TBPULlZzdK+yNzzgE9BFm6sIS/
sTHjvEzNyP+FRxiUZrTT6e/VGSYlm7CJ4d2HpuuF/hAm3pzD0y7m50zpJsMwVqGHyTfE22lJKekr
PsStn+BFe19OuD4Fqk5+F3LqZN6ZrnWxkpNWw+607PwtwK2CWzXaqR8Y9Ke5ITV8p3MwAQv3eB/W
b9kJJ265wvuRMIg4gyesAvZq+yLtQIy7as7bL7Ai7y9QIobJNdYWjutzheixRgrpaMwVCnnGefZW
UTzEtId0GhKkCqLcMK0jvSCopsKtzYUUlQUxVq/42z1ubZqF0V+RUXSpEEpL2RHVliGB9rL5ynJ2
chfI58qTFLbvEG6ratQii6lXQEEi2PVh29tvuD9dh8Qv1GARRdSN0zmMWpTFl2NVpgyP/ZDJ8NUN
ho6rxNCWIadlJxl5+bMwELe+zONXiJwE52jZFl289KMOWs9UHiosxbj7bckRTVrf1xmTloPQ5M37
wscvSGfqLBXIMzo+uvFKpFfBxfmoVgrndfrDcIdR9xc/L3Xw7WKgYBNpC5VQg6FCOaMX4s3baNun
e89I+CnhPXSBy5ZtJfocHPaFeieuu+3KWvFgDD9uGfax8gFuu2kM6uOQabv0rr/SheURH8/9e0aI
CAKlK6u8VHyIMZz3qwaV+wVW/tjpHJxf+KSSKTBeQupjK7Qx/LDPkMBDOOurJ42w1KVPxNcP2s19
rkzoVcHA8ZQrmTQZdQFBsKF0MuWDr4rqr/gAwxzc6yqR4SpOGvRag8KZKQy44TZlINkxYvsMMEw8
9EWrj/+ZmdNjGXkpLntMLnDOi++U2+MNvvhDKSLgkS8UelvMWOEgoR8ddIZvJXScm3/U4ARDVswW
XDxJzTxcH8Krfjrkel8QqCzXnc8qq9lMDoOWQ7eMPPN1KwRfUxY9E6o+yPfB4grp6bZVA3c69N/f
y3HvZGb8S5Pwz+odqMs2uubXlgLfAKzIL+LP88qhudOYPZqG8QZRN92trsYC2aRqjs2fz0rTAQ3n
d6E0ZBVeMe96M2cPscd1Of8l/M7dhx9Se6OMTw1fwUuOn2+w8xjAljHxL8+v/5uRQcwIVWQ3aPY8
uvzmFRoz2dsFG68N717l2b6/bkbIoilkojhVSLT83sl8nQh7yC9IKRcKdsf1q9KjRYbYGlDgqK6l
ORGo5W5Y3hIv/Q8LhB1CNyATHkblV9opTB2C1tPINKT5W3Qa9N7f9hzH3Sl5gkHAoNGc6yXMnoUk
Uc8nd9Z5hX7xxj8MEH6nq9Y9HfAiYfxxwWEkXDKI0vgzURufbfjXCsq4pVzMRDUPKq4U/gtLwmRv
Qo0rBMtcptlEunsmp4HPwdJ+ekY6tMom/PtVks7bC/XL453L+jQ2DrEICNuSUfQ0q10Orq9EIC4a
vAh0/m/laBJV46d0P4uLnQsjK5wcgP8fmDAHjEutsnzC+kIeB1SOb68TR839J2nQ6VHkGkfzTuri
KWQx9pnv7/KjfEepYsCq0HnDmW7puVA3M8XADRRD/zD6cb8bNw6yUcS7m7PVyBDWDUPCohn6Kdvo
B3o4dmShMFNHMP+Pfq6xZibzy8QxzvhXHyLFEoh+R4W/iIW7ussFsCSLWaxmMSJxbkrnwmGZShNY
CkKVfrWVDRrdzg3/jDIiyaTRvFMZ+ua5LtfvSrRo4xmm1INMqxiFV8p+a5sj7w6ICuZ07EzRE+xW
dZWYYakT9w9lbkrkSFSLBvzsXxaZRNNK5yv0HSM4D1z1T+sPGNFUCvtuRrblaeO2k08IPccZ4Qnq
3TTok2/SnznCxmj0A2bX7AO1EgW9Ei327YMVDbIT//W/BTFIx0sWZXvqHbNa1vU5Ow65Ps391Bi4
JTe/+UIU77tshYGLliCFwb1MRd8fguLkCIVTwx+vCQUzCVHHpkMj6ir4CGuWyQMpSZyUJZDOEkeS
wlpN0tkaUC0lwyZcukLA6RtaEv092Pt1hVpRhEqmkAAE1bxKK7nOIB5pyqPWJrwDx/DXpmOYHRAw
ZqMvbTgwYCwisuan9jSBiFS3Qp0DPZ4NPdv/dxnNvAQzHW6wv02C6VDd0+BIvEVV7XNmbKGAagiu
YCVYn8utypmH2r9nHnfNfv1/ArhcotViHbCuhyGBfVxKcJBxFfYApOdP5qF4/BmIQ1aYqqCaZDOl
ARt2oJ3agimcPQYD+3hcxDFWsydTqxUB7dGF7Z1mhYDKJiPAYniX0PTsk88hQgX5VcyYeZysjSuc
UI9MAt5ayMaBk4hiVFLPU8tmg+cPloFrlaW4bvwLaYCFuE4PhL2nYUmynODDvKh8ANcfM8f4Bx0a
OxsdLrg+5k37Tv9nczblJwV2mAI5Vt1ohwHNwXv6In81VaywmbzwzZ+MAbba2OA55TwXBJio8tah
iPM3TQG86ZnPoev8Az/Z0qmngyFHITJPoSCzMa9XWkef2Xa+97OoNXIdJe+F9LTLz/lACzJ7a6JE
toO58g3rC0lhqy9/8/S/j5HiCbiSQkM6SNSBxqNO/v5Sb1muWx5pPCkmGRWWKy9ZrFoysoe73lSD
PfJ8V1zV+3H4AKez5A5qWuBwq9IDz/vb1fuxXDsV20I27UzL+JjU+nccy8m37EBCltfjQnstUb9G
L95j0TcQcNfur+3kcKlZuRpT2/FUB2J0rAv8Qz0cadw4hOgqvpUK2mAsPQ2dYM1IJaJl704Cg+4/
YXDelebWguUM5zLNKQo1dVAFGDllvSyZRAL+ETeJTIBJ8XRMjZ2MkxSRk1Hw3FB1Rkrz/C9Q6f+V
5yZwhTT1TEWeQFx6N5xCEaXSfC10M5vno6Vm+m/QvIuUTGyL3GoqUDVHvDU13viPxhFJoeGCgZ3w
QQ3zldnn6x4VBNsfjpquDduGI3s4rEdFqohCTpn2MO48LpKTp+XbRN1ifZvIAsPq7Qz8iMk4VRJ8
+gqVfqRX3aWoJFgfzrWhuGbFzb2bsi5s+bNJ6qtIxQS0KzEHik2/E3imwF/gwvslKoRcz2v/i1TI
em/Fq1v14ijCOvzcKoFPiXOtipaiyCaQbB+Wjf2CPf5xFqmDosH4TdF+vjUa2uxU+ZYMoT6u9EVg
7U/wiOep41Pyr2XcUUyNtgO73xikz2LXPMdoIfYV2LnfKVZi7wiSbgMv5wu3iZY9AmTHTWxKr73i
8sjurrGKstnZV1xZyXV4EwFZ4/3RNawPgN227jr3J41QbZjQjv4IpgrfYFrGsRGhEnwzJ/ffu0EI
p+v0o76HRIw/QzQtwxXeWf+EFQEKMdoua+Y45eUlF2GiqUtf2lQG7WEqRAYOdRQJ2z+FtaNEN5g1
bijH+An1LZGdWXMPtJRPr9UrGAxxx+soiFkGWj2V00dyylQPZnc9r4kHsG95rwt+fDtvEOV108iX
SqGdhvfT4AT7y8aA5AsOzCWry/1JHauUlBpWBWDpN9LKjuLVZkdZh+Qst/JvPa8QyreYF9QYjF9M
2KPUdG9TUhGo/pmfrGV8itAPRkFxnoY7/73/bJna7NV8wecI/TyftHeHgGnina62Li8vXh0MzYNr
nR92G8P9vIFbGdxi9bWctnaowHRdEWyr4RiVoi40yHOyV+qjXlfTkyJOv8OiTVRSCCxT3sV8279K
tuCxWtpjETMXHSt4a5Md/UHf8s64qzOPIUslXYZii+Cn2qVVFS8VQtegfphFABsc4OviD+bRPSQB
8gvuTpS6RYTqE1NHDL4IHoybD2wH2AlT6do/HrWfeizVxzL3K/YySzKGHDPtkek3dy2nvPi8O3sk
HAnBTUKDjUvfsB+oy5baGKME19H9YBBuc0mL7iynZC8K6bRmv2nkIWeGyA6u1RkW6Y8Eqxkp4euC
KfurKgP/DQmd/BbsasX7VQP3lBwocLj3KbFS9sHnSgWN1MJzOq/NKMi59gnz4r0Ace56RjHEVA35
d/e2NHe+jN4RzKplqJLX4UCwZkaSMHkEwONbUVxap8Db6wQQX58hbHPU2Yq6sou68X3aZaD9RpUj
y1WERC6j47PgWs6LxEyfQLRvRd5N4M8S3fk6pvKhWnsvg4ALysApswWHfx971uYH+0Fw1wZ3gEzr
fZWxnhwKvPcL9tTwIVjHOoEtOSqQ6NplQIrVKsFviUz/ZKcNlUuNSo7iX4LUeYoOv7W1nYM4E0UD
qYt/vsee0wS65RULuPXkcZRAz1P8TI1S2byw7bEGPkz8q6QGJedJWh/NB5FCJe90u0fHXdQGEf6C
Fu+3zyNS/SalLT2+4nh3qTC6K81VnIJXBzFmNkhP2J+uTBChrKsGyS/IFelo0MnmieSkiteRMhdL
LPDlblu44i5tHbtEBwEg94hXvIEZvJhOOIuwzh8DwvDmMZsePMGchJV+hXBetZpNfTbmvyzBnIWk
5ab3XjBI7KDdcviX6iAPAsULGNWgc3rMx1Tq8BGA0NdhKFwFGmkoezbHvEcse39w1MxE9mgLHucl
hE2pDqc/xlw2VoclG8cWrcb7WWYvJUZeAoeYdLjBG//CP8Br6VrQ07Mv+yikflLbCWUn3RAKmmHv
7gU5X8trKIQOVfSoBGfwdXl8Clb9+AUhjOBm9FeU+05dPRE19YkIzNq+jFd8BYLHlcpAuxknFrZJ
IbzE6kuv1LgjIBDJssT72vslP9yQC/8eD34U9MWtWv7n6TwkTUiH4mDnaYwLXFWQVYRrxb4HqfaZ
tUwVUXwK2ugLp2MNFtNUN1BMeVgnshnXLRrDF3/WKiPmFM4E7qVrP23/YUl5EE6LviUkYQf1ZsnH
qKNM6bmkOQcSuCfFv3ktuG0oRpYuCGH6y2fwx7fUjiHNRGKUT/Rj+p2DhNvRm/ni3AMJxc8au3Hs
e1GK8lW5juA0YaYExKY2bR1X9t7AlqJEeP7vlKpuSxnaAuhs5RxEm9E61IAboruHDHRrJUqWiBPc
0QQ9hXd9WzEyCvnBrrzpQfptJB63zt5ALnZ7t0l9WpXamMhlCmqOYS0ysWF8c2+pGcVZ5NI4e4Y0
21RSqRfpYPbB0XeoVnEqyH5fLQmWj98TO6Z7koij7UOal3E2B00zEzcExzQDdX3o7R97LT6rjVGk
ZfE2tsm+As5qz5shhd083e+6bsQkoqPWzi1FPPTa2jPDXMo1P+LWvkrliNp3CQa49V2xSrbccU8Y
I8Q1kkDN2J7jbcIVPxzk0I5CIvvBRpRywMQCA9E/Eoi5yhGHx+8ntvAnwsYOQKCU42PO5Y+sRia/
psSlA0gfL5DjwqmBlKL7hyOz7a1hr2GPRc7xzNk2GnLw8f8EFIdTLfPa4sskfLohqhUr7lU+koq6
1WNQBVy3VcenUhWBO5ejLhYu6qe6kfYHC3wNdn9hDu+K6zRPElZgEgN45Fu11f9YeMRqUxCbDzAK
Zbob9n8RFMxfBnokAfAFDqvfNJSyduq9kLGxgyVa3IkERba9OPX2grU25xAejPMuEyTs5D4fbLMs
nOhlj519bj8NPxB9T62MHrW3JhqTobWinOF2wRAhGwk6JvnPOARqVqAxr7shmxh+jqS5JgTLFUR7
HxJvL1Q8P4QV4sNUr0uT3VN1hPoQC24Cwd4h2n9iSbE9iUumE54WxNtj3e9dK7fRz/Vsv3xRfoPb
Thj8FHQOXplBbNiUNgOfjfI7W0fT+6kY7ww1MdLcXpZ9o0Ca46Z8RzIcwKaQQMtqJmlcOPI35hpb
1SDz7SD9MbzQu02ilISo18MPMJms7Lgj5RofOORl3StEo8vvwOAIF+vm8KpS8ZiRLxgKXLdACzxC
sjguiIv/lEvzin75uVu+FnKmnzAXk34hKQ55RC4dM+895o4JYT0HGAwak3XCbA1CNyZro2dxtinQ
uZVb93dDXCNrVRQAokLg/WeihWj8Jh0fDRDKARpI15MTvtHTSgPc+6I8VR1uAMyuuJ4hYlm2dXJ1
Ms0a9YFhZLCglHMxqegsPm/I8DLN643y3A8T6SkOSbuR3SxHB0ECvJl/p5DO9/8n6bi6yNGW4wyM
00PxXVy/1BmO3nSQhRwiU3teYsQnfaydqnqX5GwoxVrspprk+LFBs1I17dX8/+1YJWF2eqmh8HIb
PTPzn8Z1SQRVB7RqiFeseRRTzkm4s9OkiWv+NclOY4DcQj/6VV+UIpcmohCBKcsP3JCXO9G/6gZn
hiUPlSIq69qO2/t90xoDzs2hgUZ9H4Knv/TlNzpzmPOc3J5VIqGL9Do3oFWUGj4G0Xe3y7Jl3Urf
PdvPvGlPgwRGvghs7oUHCk29BgKUwkRLPYJh8j5OKiVXnV7RBXyHN22E5NhvZY1seElCFSFUfFhQ
kcQbcdr096fTcPPNxbFM+tzIipvlF2H+PWxCu//V4nG9ErljJuQfnRt0WaO+eO0RXpsaSlNnWW7Y
EukaPtoojt/wnP+4Boum+crQXE+CxqkkT8VxxzkiW1kE5lNZXlQwIrlV3LJxzgJZpqKHcmSkdHHn
RRDxdQ+jrkTMcMn2UL1VjSmu2/JXy0YzcmiY9ucwMhTVDio/WDXRGFL93YvnfMH+VlYCNoH3hdoh
NvitF62Y87qCeqWsNLbHjJYC5dlt9H6cSaQJkLrd6EtCEszPD3n3gw36HtZ7lZlnq0kBy56h7kOV
rmTqq6t9uDUZ760XeHvDLBFeNO1EtAymB4NE3QGr+Dm7wTzyfeXs1IDxq8xMuyt74v4+HQmHdnHD
VWr1alQG/prjn0TlPKIwQBlgIQo9pJzS9qw7Q1sRAt9MLHTK4KDqy6IVmN2LKTQNBKFerZn8clTe
qbOVjS8t0/0LdLlYevjNqlOqkMsyn4n63DxnT0Wya+3ZunMQmIKHJnCWVun8vD+2I7d9zzkvvk3X
bTCFVyQBGrQaeSN0oVOW5Nl6zDAYTlGq7DAstz8bqUTqU5lcNPwPY4b2TIMJPQBgMeCER8ZYUkgW
6yzP8Wv80/Q8j1T/1PO8tKcspMQSzc5TtED+gJWf8BRIMVlmHi1LDbnMEc8/UMFFIXJfmxa0UdNw
1CjtAvfgkL/3t8RxX7vqpUUitVqZFzv7D93mmAKYNFZQU5hDmVOptWMmXlbYQRPu01hDPkMJxBx8
08TXeO+7Cc0zVODQ0U2ZhvFVZ+8/5WwVZuMojWlWlR711m5m/+tYB7VKrR/6XdjRrcVFP43Pjarj
wcbHuyE7SDsrKtKQ8MBj5Ok5LLWJk9nS0U8lCCeqLc0OrMU2yWaltjgYq85vPAvfokfY+/GyBaMv
OlICmqY+5Jky2yfOYiANcanpn99TVmqeW+T4RDR7WGPK1m69KFNv1nkNNm7zaRILXfP4N1yOHPyT
a0EdWuIj5Vhfg1oL53ELoVDmdhmUfXiENLm/Qin24P1Kn0ZvVhyGxN9j8FRUc693ZrY/6zxvzyUA
qX4QBBd3eyDlNaoOyiM1q7DAsTAU0eSOTN4If6gc0mZTaRFDVEoFFi8Sf4UE7GPm+7jMVx5aM+Qr
KaemfBLxV0avqUlGPxhRZ7H9DUwZSWcGRCqqleEwlhUE4z4yHOeHixIbF7rqblQsW+p+SWbbqlwD
tQKKM0c7J78w46v/igv8dXXFg/Z9Gd1KZPmR98xX0XMSyhuCWO3xFLBypDlsDrGs15QFnF9yyQM3
b2uhODvDt2SQjs7hzWKTvV+TsffsyPpHRgJaA3WeaaqcS/vLAsajUyoL/qSAEUhRQxqpsyUjKY61
VkB9fogqGtSJ/6sc/Hrx8NZghv/Vmt43GdeusLIJNj1tJiBWGPC6NI7tYEJ7/Xv/k+AYjGerpoTP
BOy1r81nzRITK0DgdRvK7z7yid2DFF59yXCqBOzcueqAfteelJNPrIPFOhNU0nBIf9ZplHHGiB1G
xzynlDetYflStRPmtypeutU7g2rw8jr1Gs2aOGeGUKnG8C/E1UDdy3fxGI77rmO8wD8sq/9GAK+z
oTIMXnxKp7a6Baja23qNLly3cd3KBTib4zjKKbcVp68CeItUPQyw2wSp+OJjmEV+prUFQLV5oVUR
Hz8iQFM+yh8pCW4GQ4RuBkS8udQnYNIyGEJHifMmsr4FJNaBtNSIruFFv0vEQMZQnedR6nY4WySV
hUaZRSkmrNJFKJJE2UkhXIXJ1ekCvwQ6uoYdEwcfvxcLHrUhpyEaqhQni4XIgbAmGczyjprzx/Tl
s8EMFgtGUfn/5RbSwk5pRwI9c5No/tSLuYuMW26VkiPdRpOy75WpoZXrPBnhY+Db2aCIVCI1pBnU
wJG9uHg62oPxIn7PDTRiYOD849Gw7PY68c06M2DhMTBnZbJ3jwGl2u2LJnVm18KrfKIxl2oqcW1e
XkgtoLqTg+gGlYP55RdTZV/3viRwYzrPXZIZx2Vxs+RO9UAYXykxPLhNl/ukt1gj6EYUe65fJKd/
/DZFi+lve8u49LQQ3381HGKYZ8P1kZ02c7sUeEeI9afe6BHL78WnHCmYGDSeF4YVdDgtiKa4dqbH
5k413GToYl/1HFJ+rkjpGfy1WHpnUSX7nquK12kwOtsPFsw+X+pjC9dVPXvit/0lHf2cnnXbLVMl
gYqdJQaYDhjgFNA+5j0QL3JAbzpzlVhNutjFxL59aGp+vzCoc2NPoQVJiw3zuv2WpvlVQOAgTGVG
t3g++bQURTBg2RNsPs6UnJdMsRvRrqolYoFhEb5SagaF1+EzWUB3E12f4WxEzf0CbEXoNlaa3nFm
0W0MGrPA5RxjD8iNiTYWwP/9s7BXo/b5UV4nJRqXDxHztJ33Kb0UNTDru9+2RTvJJ9Pm4OOV69yC
jwCJlS/fKqvCF7vpNMKpK7vrkBrIJolxsF5cXdt/UVrTp+fFI7Vy+3S51BFUop62XhEVOHINezqx
2SXuZ9kJAcjtD2Mtu6eamjSdSnXuEe4/ZZLzrACb5yTwA8f1jyWh1nHSmwjhVce6sSLfJBCUxyqb
BEhOhzFLc8nT2VU2T2UguFl5XFSCd26e5xWItgGp/5vvjt3sEn1KtmCgvYyojizqDSfEuST6JuOg
PQK8QPfqcM7u9NzWxacGl0BOO+gd32PVgzDShy9l8xbBSp75Bnyh/W/Zf4Rz1uuW7xH8B/11EfCV
bFzuLJfY3kbN8mfY/7ceKGOZUXk46UXjDiJRIuSzzeds8K146I5rZbzl+VuBF9IuW9cOIZrruZ1p
/un/B8+ilkPrOYr01TSB9XQ1O5YYHJRPV/HRVaJQc9X8qld8aumOokS9TNjXm13QrOn2Nkom8JIf
HHD1HWg0nu0FGTaDEa+KNER53j6mwiVGUKz4jJep7K+37LsiiPOKK2ZBmowNlFTJbQ0uapXgakBM
IK7fUgtc+v/iz0IT3ycPYJ5Ap8+CeZ5Q/IJWWwoRV2OUS7dXLWbhXy0Ef/r7LkAIfFlEnV0Gqv/F
cvqWZnd3r9ul3d6aqLRZ3CnF0opQkqQLMaCuWQ4zh9tTqpM18uzQNSygmpDgUo/PeGou0Pv8UYzb
WEK4OdEuBRrwTG3GxGDzwfCjJXl40xGk2QAaJH2oIUG5sneu0besbg4OwtJOOzx5RpDrVGQ8bz7d
ozyLcDDEIhTn3ZxDLIR6f1hpctMmDnQtLVZAHmKKKalLaLZEpOfNJ6j0o8j97TWTRQc4qS4BD1Qw
7vMhSlh6/ec18n5asPUp2L7tshd14vsZszqGjbXxfaY/T5xDzgvPQqsnHDWctTjCq4CERirf4z+9
OobMk04wZC2bE01HuzGqupQU5Q9fznQlykruw2uD7Ed7c+McpUTeYR9dKS6Mj6fLO7MkNUK1MZoB
VzLIq6mTaAYtr7wFmfF+M271r61lYTb/BMI4/s9LVAyF6xD08HQvk5InzMDQsB1Zmt2NyJXNqpSb
hliI1aom7UD7ygfvuHQ85V71CZqfdHzL6tWqfDANkDbW4KoepY2nM+KMSfcWixHi9t5Zi1cauO2E
/+lWURj/xJZNsxh32wE8hmm2YntNVZR0ZpDY9SqlgJxIAdV86cEZ2n3bZ1TIdii9OTWfV4zDyCtR
MraT9JqkWJVUSCbRf5NZvTpJtsDqbhGjGDZrfpqQq2b9nMQOEX3usDh+AviPdXcZcvb9lLFW2MXi
Lmw3YSkfH7cO22nGzxaS3GVJLLxYv6k/4OaJyCH144cxLz9h2x79k+5FKh9fhofQU2I+82N2R/jE
hrG6ujQpV6TH1pl0Tz4BPnxxSUJdiFvq3NYjh8B1kJHrk2tnSuKd233bPCsrBqnPG0/biMnrOYE6
GL80/mMI4DLCUbATkN/BZg5X9O0F+QqZs3e0H6lMVRLgRiy+pyOfZuhlSZM77iy77OdwJmG0gmDO
3YxqkanwLHwqQQ14fW0/vWGTjuZFRQcAQJo+eEU6zjbM8cU88BqzrTzGH15x63kCLXz7smoFNYe4
OemJ7VNS/XiBg178P92/2PL4CWnkDWOs2+HmL51g0+TXBnlCjJlx8L1dqTN1C3vESe/FMw8Gkq8d
VQgl+JYKljfPgJv5l9Ck0vpHUfredKVIGxSS10qm+NkcFGt4zKw3PZPGcuYaYdEQIeqJjY/uw6ez
PuT/0VOR6sNSx54FFW21L76kz2NThvwzy4HbHaTVz0WFwWq8Dg9tCsjGNNxQsvT6c6DwrTWbDz8d
/xnsVK7C0eHtOYLXzSem9vyNEi8nkJ0Qu5ZlyYCCL20CvnO/In9yvwFEu06Uhdu+5F0uhyxx0MkO
PcwBKpHHQrdNS9SVkOvlLql3l2ZabtDrNRLm8oJjHHk3Q6YdNtvgbW4b7m6jMg35+MVhB9Uorthy
yWGSRUk5P7lGspTnIfQaE8phtnO5jVGJn+2wyP7c0JnDwkkKlekSX1tBRnJNtE9EKJtvntHfu3U+
L7+Za7s+dIXt3kUbVgnJ+I3WW1A7ku0jd2HeNm4WPdQjW6D3PG+ift/FVtQhYkJYTkR40tKbj4yb
N0VRDWDXnTCMFIqKvUmROSGH0SLofkxtAl0fuUbTILtp16Ga/cvjGBRdnrNYWq1I+xWynY9Tm7DY
TmEhA8UhmxiQUzSbW5+uALT41MheNzbJG3p3pqzvzD7Dalm+mIa0peGcdL4YodYLSXOGwbln0MB3
yniv3IqR7lfBAWSF1o8AiGSAPQaJm8pdl+Xhd+OjgQI6BITms8PP5M7T/gSRyfl+OZfQzmHnroTX
bJogq55CpnFcEvj7HglysbeunRNIQBjyuzzvWWv1Hzd9SLzKt20ylBdOdoCODbBVurZmU6hldHAp
XodnsA/iLjSO/y5PFhlYZKMmll+zcKXUEnso0MskuC1XQtmeAZr3hORTBQ/pLI06oBLYWNFrZIIA
G6QCB2KdrUuDrgYAPLyFq+GNeirGmzIA/igPxu6sLwwXhXiI/BPzfZ89rdZIz9h3cpHT1B1Xprs3
ZsW3dMbLwtlb/7apHroURFxJB+EVD93AHn9KucMyKbQfX1VXFxXlHwtIb6eRYYPn3sZNrafXShp9
1j1JlK96iW7fLusOHQxIi+17wTbCSMkiriUOS/kidvrjzmdwPntdXbSr/+2Ti1GQiLeSqo0khUGh
ABImTJaCVmbSDgYHfSHXKG0CpMrSmeHtBkJAFnijm4RZERr4qtmuKGBUJnTfDx9dGYVehG4PXZAu
0cBPyryTGnLZ1UdTwl7uiCjL2xHG3bbw59ryPUvfMQKXIy5OAgecdoAJWnfw7PB9UYuqDloz+Dcv
ljZ0AuLKntMfvEEZ2YC9lw9uo9fY6l9hepH2gaRGEdxb6srCNj8hWqfLjEx3NQWA76t8578c2mMR
ohBgPy6rcucQZGoD5T6bGqrfT0eCWf8qPy2UlVkHM0OAbI9jU8CAHYH5668Z6pmy6giqoYNxFNr1
yzij993R3MoTvCJ695up836CwmI8BynxbIfsX2HVCoSe/7XPfz8oQI9NHjpE8l4LTTxs4FzsNFOx
NTmbVqVJDLEUz6y1WLVfho4D4VrIs8Iy5rzK9pxLoT95all00MvQEYiByVBLGWphOSmw3QkawBbN
DXtvgIjIRIQqBWdtgQbZzDZc7f4a4QeqD8KjCsQ3+2+4QUuhYq/LeooMbRCVPsXgV2uWgF0JWQPg
jO0WV2c7eLxLSBOafCPYEFuB7l5vBV/3ZpNHxq7jCBpW2G6MnKxO7E2gD0Nq1D6vk87kzpUaDqWK
Elbpmg7jWLKjHVQ694A7fpMnPugDsrU3rqQ2zHkNy6LTZjMTLKNfCNsWY4I6rwH67ZTmdxpgVoVJ
lwmJTYt9Y0sEhAZ9Vl6GRXP9Qtgi6ENsmX37Bt7GfvnLRmNlGs8huzSniIEis7N+bU2ApcTZu+fr
IOVRhnzKR16kUpv8MtWuIX7x2J25Awqq6Qj316YdThDz8t3m/KfU3cVa7TYM901pQORFXFRfzKQH
sJS6xEBrIEr0feA2onGxwnJujsVXNyYq2oI8G7pZeaHSOIt7Y0w55yNpZB01hz3rjZ2/dVYrDTad
zY69xMtFvk3NjFGWyyiDbnyzFgF4G3OrGuwMyC0+jWi4FT4OhKuVby263BoXKED1zT3rne60MpPE
5dn/ifPkfBwG18FEVB7Zk+B6tb2NbW9SlE40qSa8G0LTQY77eLPg9q62YL+hsahMCyA++Ps9l5FX
TiJCZTupbeLr0eDiziKpGPEth3kus5/qx7c54kB+CzHCBrF/h/FBrkkyQUnKvEQNgE8CTwFkUMgy
j7ZloIKeLhD/jXAXqYysrCVyxsS7E9hhFdXoNo63RIle9rlWVDegb3mWYgDRSPWx4XEYwGbJtT+m
ngOyaMi/4Jnfk6QZgUaaMF6otlTxdWK1ww0m4SzLvUtQwDqKDXQF/haxXxW5P/m3Xn2prbPCVYT0
cp6fXVl80dwcxZj9F0FHA3/9X5AamOO1yVx8CYuvRZplFjqFGePIVqS6dWND0319v4vZXdVt9JxP
I5/Vjygm5vlH5XoAVlt7ATHVGxFbRLO6wT5/9gzQpiGTYl7ihjsc09HrqbH1MbGBK5U4gURqX7Dv
1hOgDbMt6eqzrFHb0MFEl3yLfhAO5KRqJtc3w/IdOGRU9DvK+wziTWwJm344uepFrHtUsA4HWE4h
upiKs9trLf0HpG5e6Lavg/a1I3Go8u8m85QZIiIeRs8K8GmUZ6vWHdMn1OWSuK5iDuC92mDiCOau
cVIYLLgGchlED8G474oj1WZyC8AeChnsc0GP9cznC6xrmJ+mVhdAY+DMnB1OXaz4oVP5Cv4kWhA8
D39TwG/VIY/4GKp+qVgwipoeLowD9Q3MeNcKWDsrmPdLAvN0yjlSpvXfbmOYW+rh+o333ylSEmgu
6s7J0rrahJ4oT+v177rBTNlhIgkT8PeEkxGzW34W+Qy62hNS3B32qNeE7JJ+R4wnY+PZaeJdhVv6
FSshjegASaJX1/Zs9Em854xjqD9bMe1quZHDS3dWgQ3iev7inApwauu2QGIsdN4DhOPftXzcCEay
2CzwdERgncNurQXICoYyyL9EbURTpiVz4YwCmTesZUwahNTRlyhDgrpkjYXygAvvzEt6NCHJRKdO
N80qsfQKMWXmWcLQT9n27KTa0YhhMvpLWfkWqwWTUd9A4cVOWQW/j60HpTqL5pBSAVwhdfruiSDy
lRgGPaQ2RJW/vfnAyX+4oWCCz/+fcIhpX0uww0TXFksMoqfF8Sxgt1/8qRpBt1f/qXwH++rIilJ+
u9NrgtuJt24bbduMR5AMApsF7jvXPDPGw04BjhlLgTTOhy0ONGDRK8dplmsowZAYPMCJm/60sbYX
5/v6s8CEylL0/Myca0WC/jOuA1OVzvFAJZhl9RiwLHXnfpDKMOGiV0H+GQAV8M5iYuBRdF5dnuMW
M9r46QOWvLoZl3+5NMVTwI5ieFvXv/W+TXt6Dfe+FSA0wMYLxmHS+LZvaJLqKuO3d89UUcP1FOcH
hZQLfoQQvc/NEuWjnjedHDjNHVepxr7VHOeJi71QaU/Nh3VntnowehhgGS3y5xreH2ETtcK6i4Yp
ZCrnOd4nz3IqvxpvfOwcbPS8sALehh4R94dhlpn//Ke9BcWEpM5TPJqYCHgbeuFfaI94omt+QK89
8wJcufa62Gzvvf0NpubN1+fD7xcK4axKTXA0xnbLW4jBEQhpc0faubpbufIFHpXsgMdNYoDp+7+Z
IQGuQVKhczXO7UGUm05PEhe5+7iJIbsgo/nAOvkz3E3xevJpBSLmYuPA5ODC44ajDO7ZkbVYlPd0
A1CieBWZrrJqQJvidkQ584Lq2NkXR8FnRMF1eSfxdiQzEyUIV6Wb8pFAfgAM+UZy2bepf7snMyf/
FgwraL0PVF0jzIaiXm0YHZ2XUlX3s2XD20RjYPFsyhn4uxKgMmxBgAT4nceKxtsCb2/a5XdrcvyF
KyzT/6UB9lXFzeY1TugkHNXnMvQb/6qvmg0M+m1ImVRcgG67rfqfcOv0+2PblBr7+EmqT6kK31wB
mMcKiAFifOVz2hwvUW8IWi3v3wl1wuc/+cIhsK0tGrWOF1YNRS47n6fi5NK6DPFNPziCPw4p4xUv
ZgIJ7bFlYCdrLX5kjiR4VtC+qcNN6+dJIGp7wPq0wRq6hnQqpTLSsayr7ed/suN0mJYNtT4FWdfv
ukLV8NtnozhtGvWzepMvsqU9GwW0R6Li8+ugDtoRRq7ahRuB0eyd6iS7T1TnLksDkQz6fzQa3xkL
TPlrSyB047SqEAyiAnaRmMBU85rfIozZZXfZnul7vZiDZY/o1ER2d9Lp+hrolxLsQYwCore69VdD
jlvO7KB805nbh2ImvIj73EOEj9e790CZx9iAbuL6js7uvNUJ2oFcV5WRMbkmtDg63pr0fT7VzYnA
GCzq022YIwNKXaJBFlyKMSTpmFW1pW6bCqX28fAVrKO4S76zB9z7ZbFUu1pDx/8N45HNmpS4omhA
ZqQGKmqWsYxio4hRNuSmcEcSYhmGJAy8ZAz2RXlX4liGT4XPsFfEaKVIg0svQgZQKeP1RHkeP3v/
II8IKSVmhrzyErRnM3vXewU0HEJT6okIaE5EpNW+MvK5HK2J5GVlc+LupU+an2osq/UyFHAqL273
BjqweWaUeGb98GXzynh3FGc3XLMlsCe0/9RF2EHA9485eUlSosHMAvZHK536pd4RVN0AaMmvuXXY
2lOrwaUYprcD5HVDZkvZ8RXy1YJQiuIPxJr0L9adVpmudb085BnzY8RTwn3OJW+89rvH1UhdoFEz
FQiv+k5kIJMc/XrV60yJBRBDwGP8rFvFG7o55Q05coR9DhnZZGuXi1iMJCTtluR+X5iL3/cSc7pH
qhRiHsxveY96x3lvsbCAqUwYNx0f/Aag6VY1sc13SSX3cd0XKioYOEB+JY9Jw6D8zAK6iwAM279w
5ylyYht5+hyqnIi2g/hB5FegGn8HHBmHoDSeYz9aCeU/IcU758nlmL2rPIJSV/zWw9TClj7iz8tr
ikvZN2755AD1lKrS8SLRXXgiH9AsE9XrBiYKrM2kuTSr8Z/lyqLRLawWJH9roTOTa6Eq+ZYOq15c
NVBVwZHWwUhsVrw5qHr7GYWlzoPOc5U/UUPyAxnZu0VX1ItLJsMDPepB1DfYFUdQbqOvpGsNq2TC
T2Adz7uimh57mGSp8xXR53/Wwur4G+0/KBsnauXKla8GYSRVrKexawhDaBxYy7afIo1CGXfh1oRH
BnjZjvUEUCa0Qg6cgtiX7M1n7Y9CqYVKNUBwTpiqwOGSXClcV3yRckZby90RtVgoooGIu2VAsLLx
XsgwgrCnA/IIiXr/Nl64BdgKGO90Bw2ZyOLC8tayQfBFsETl56tkwFAEKy5HkttIxoWwst42y/c2
dLKkyAQ+o/1vk6gk0iq0sPdBHH+IJoo0d+4oGvn0eLvjCu9Fe3MCfsR2ecNOMYF9y1yUwGotiH09
32qpO/PneMPi1PWxnIsX1NqNtc16maioy7OtLGVO9GJRLO8xj2KTkFKDokfUPjpZgvXlERz/okGS
ku5i3iFCmiKlu4Ji5Z9kaf1g7m8InxTKUtqTVyVs99hlBxUSa3t1CYDoYJnM+GBcofVu1KDn3Qat
220jtVdrJQCjVNtSlr5jh5FLS5rj1FroGjjS8AmdLwFYfoIQ/nlmMTSPx21kyUgpPRzvgC2i+nCb
w+JcePBJbsaOP9CIxfqKWH3aAF0pIFhMJywoEX8KcY72zxHVwOePA8e9eBcKuWsoSumE5QEKaQES
TRr0G95AFxUBSSGxUTCBCpPs+0sSOMMG8Ghb6TaULxwGr66zFvtyCGmC+bco+VsFQ8qGKt7G7wQR
ZkDoDDvSBMzu3MCQQOpoRvJZIONdG3DKVXlJ99bxV3UMQm6uRosaDFtQLxzQj8p9k97z4GdYbPa1
+9c6qvZUA/Z75nLk1DRrsvxoDQBV6N8PDTc5QfaS++qfi4AW3d/Q3FMPcdKW7lZ9hu1lHbgFWMwG
nEknCgW5QnSO8uwqTrJyUL5neuV9nr6nRaD0rbzRQxrVslNXvcfmm39MmlcG5LySyuiLHGiKLxP/
lPPnshxJV9pn5F/kyWUvvhyMmqGp4Pqy34fMQGNFCcrHziV1kyz8/anxCuCZ12QMkXcj/IbwXxG2
AFkCxL61+O2a90CewlBVu7VdJf5FdSK/47H+De0kMtxv/GsAQcq/ze64gpxM/lFmkdHDT1EjrpPb
K9kOW3u4V+UV0xzHw+c253vtInpZJk+sDoVpuukEo6UVk66EMQebTNnWIOwI40rIvI1SQLU0gx8j
XjyhIcq9I3hImPCu58CEfyT1j8wrgGsaBA98hRa+Av/g92lN57u65jkZcwHnPc+rOSLIu+YwIaQH
EmTrpwUeMghZNY7vaGAuSw27wc3hBxlOaVyt+V+8qsUEZ5g1fXFocjpJaLKJJovDqWQnQlkaeAGa
y2Mzmh+b213m3SSsg0QTAcvkR68Rli6eqnJM7fJMuKPHZXbcInqUWACad/4Ix5+ILDoBNUnt4kID
W1zkkA8YcxzGEvHLItSszQU6l+pBcDm8Yyr0X3UjW6WfCyiGsPcC8sbrZ3Vgr07W1uIw0Ht18D5p
iHpOzS4nBPdwKeYI3Edn35UHutx8fmIrV8kTCoIuZ+RlVJF+QWC7zIDpDi4wQxkdgIYGecP+Sl+H
22oLeIr4ge8zb/kUB/hd3WKPhVDtPlGi2Q0C3h31HG9ZZD+jeqq/Br2vNJ31LTct7sIBg0/Y7k+2
LujXJM3JvmKeE+Gd09uNAPP3hMxn1CxXAqnTe62wS1Mt/qpr9gc4+pHeMpoA39uhTgp7qbV08JwA
j2B21Hfy4menY/0w0d0yegMPc2/ELdUIz6764xd7T4wmZgudFYkn05DOkBIUUhG6M+0ZFQKmnQBB
W7YYack3BZ7axpOGtsbH/w8XsdPQG/70wla8bzj45nOJAu/Z94fCQ+XP5/G+AyZqftSpxLbNo0US
lquhcmRaMceijAfh217q6wakAT8UCRc+PpiXoqvMU6kGZ76MUbvJ0IG+C7mPtL5sXaxAu0KrjYfp
Dt6ChXs6GirBVj7hIVzxvZjmBDbvC1rbZaeZfw/SA93J3p2H6Zkn3HtiC3xzZrVZIFEupAUla3Eg
lTWjS/uWjIDcg4BVMM0txqm8WUFJdmT0g2j5Sag3An45ygOA+AvY8AhD9iqy1LQoos+FyXCv37Fh
xnomWVYvcINoxYy9kgEQB8WVDavFHb+C5QfzEyRTv3P1YBpEBi7a/l1gCyk66vI2ujC733vkluwh
397PjAWZSX11v3DkqaIgeHO+g7H+TTkDeVOB+OLnTA9ndXfHkhFYQQRiCJy/Q+zusyj7cB70qFJd
9W7dpczlUY54PML9g104O+M7ymmPzbTZepWEtcQRzqrBcZFItseEWOnK4Uvhnb+Y42f08aYmN7t+
ajFeZqh4STvJpDwtmgTSZMZtTluGX47B6DrKIT2Imsd+W5gNhJoBELBRlXpE6TP+DwzLVALqwCSm
itVsh/xpy2+pXbI1Gv3pvNDy5bHT3aIvyLE1qF2PqD57uhBfe99syNcJFfo5h6OP/LwFVes6m+PX
Djl5XIMapMOHehOrOtIUz6dHVP4LSk+Kli+CJOJH18JRPEhV563J2N0ug0sLcWriJ5IWG8tbMxU3
koQmNFUGABNRqMBVD/bxrBGQx0STgSGrq0WU8+V61vNI+j6uTRz8NXTcddhG87WqXdujQnVgtOhm
VaNzeKmn72uUS6KURYUDuG5+5FAr6xN75c2ArHbSph/z4jAfL12bW8WycYfCNTkfAFdVDSFyxQ7n
coSFHnwoBFQzi3BaVLtKHi6R+ETcSOsQGoinIXOHcqMu0dTI9X26OIN0T3lEIC79xRa6KHMC2h6F
Q/Y04OAFYc7Fanew6c89eqQrR4VLc/xnF18trkHkaGpCnfOgfXfdLKHKK01AdG74JbIv7gwMTI4B
CMj/5ugj9UJcL0JMUdavpHpER7UnUlCp/4kDaR17t4o7oIIl+djITVbgw/RPP8j9+Pk2/V8B4u+0
/sRADgoSI13YNIwvyauo5IJiMXdf0niPCXHYjfuss1mcomZG3J83p0qa06eMet/5vApD5f/NnjD4
4z1mtOFbpuJG2tDayM8ZT3Sz01JYV3VQSReTeJpnxhcBw+zXsD3dA61aW6rzppXYweXYcExjNS5H
nW9JZWFz0kTJPEwa1jPVdMy8I5iUw4yYA/xLncpyyO0wrjcCB426V+gFuqpbvOby+WF3yeJclAyI
Q9s8HnOR/ViOIMPkgjUjvoPnoiWwgAWKIL+JdCSlAdVNJ7arqxyp0X0TwjcB7cfUastncsz7xTlI
lkwr/swaCtxtwpl+1x/4boVIBY2/+DmNgnei8cQbK7nvXXkb2e86kqgFBoCWJ1zK2oc9bWQAMjL6
Erqp/Suofqe9ozS33vwznzkmag5Z+3mJqs0b5D2wt6+1g7fLpNThUGeOonEgvOQo6ERaGsabyfCR
ICNtmbDnt/H8gscbfVZzDhSI5BYpnJPNWFzXCZM43dL/BpChT1yif0l3o5SRKn2evN6glAOA64Ak
CYknlT7ZMlhMisp4sZ+P8UO848c+hMqHAwZTGBkZzied7TPTaiRMVi8lmMHjSDoz7JWCOZfM9Vbb
QJGK8Qa2ZpOaxTPEgyJJ8I4K5skkScO2s2j86dwSgazMcd4FGjd9mYvXkjifANSnyxHUWAhnL93J
B2BHUkhnBbFEifCwwl4jRAJASkqXgiD43drZpHDHcI2I2M8Jtv75bZlDGyJOfsw0S7gyjaJuujQB
QDtp+FwGYKiWot59iMQA6SGcnNMchldFrMRI5siy0k6BfGl6zdEmIj8XirJ7IZlZJOMI6Nc7bGaY
jVIbRgcFvDywvPLrMxIzIk2PTiOwJenavymnAl+ruupfT+nEitF1mEtH3yvLM4rWgIHssc2bXvJN
Z1pkwfDQJT2elz8Qq4d73ZSEBxdzsrR0amlEVw2C9w7Cgt3JDNPnIqqk/V8JTO6/l/UMBkqt/euB
nUGdQWGD2e9O2RbPh/3dvFBSIb9/qsVEAyUNc09oJLCn6j6nWmMDn4M77JRw46PuzXUN5zGo0SRN
cXa3/KeTGg4C2PXZkTwAWvezp9GDC6tkL3sbdxZPYafTklFlXMBPZUABMnJlDQROiMDXh5mNNJEn
HaW6kwK4LdDaIF+h/jaT/zGA0Iqla5VNf4tKdH+tAdgrTUX8VF5WiTC5qFNBDLiFbcyS7zwPRTli
ge0RQP8rNUg2DT93bNSCEDWPWCdgaoATSTCrCVoPCdERY1QAGGtrkmknGyKJ4/ip8oUnQb6AocTm
3p1lnwX7+ht630Cp76ajZP+WlMPeMQirhmmDrXb2e3klX0Xwrlbt4hFuGSfbr7t0kM8O56ITpYux
4188Fn0gC5S93wWEBD+iARboPTINaI2jKQ0Y54A8W+6bWbLgI/ahMtpJseN1H0trHPmsXV8LMdTy
dboln3XrFoaPHCkV+wySXuxxd/iMFlk3nTc94pR4dz8FFZzgEe5lf8smJcP3GEu7L2jqjs+pMY5T
DXJ7/eAXfCxR0+NiVPKPt+4fx7riwtw9hZXEtJ6Pup9T+lAZAOa8RjHyB8qIdBe28aexJH9jSGzr
IVClLFHy13D76BR/PHFAtewbWjayaBFY2xQ/d2/hRgUGeagobT9quWJCLA2o5VVZRFb9/snUGRWU
Yb6Q/hU935oJCvGN2Ryk57KayJcDOeKu8v1JGtWwCh1CBsP+jA5b9W/WzBfP9c3QfwMZWKi5GZBe
qqXbQvPNPcQuT0VEccAl1mHc7iZ2pfhsWRT3yXiaoNRe7uukDon1s5flgFr9tsXS3GQVm6FOCuzE
cpRmpubiVRQ2SeLJYS8gfJiE4VtiDJkVQPRDDVUUaspuK74HuDZUqvnlAQntSqtajDINNbFtK3Tu
9dZ88DcDhYFkY+SPMXpTWGxHIPJddI508i84ilnW9f66yWHpqSiWFvcnF0F/YJf+5wO5i5gmjYsq
JcC5wNWRYLxgpBT5poCmDpvPJEWXeIuKMWwQiozrVKNMD0pSMtFhM0PtKGF0jXPsWFW0oU+lxVOa
II55DkEpVr3ZtYn+sFDKAcrnDb5+z74q5uPAL2w4170MNQNJfCFD2DJzKRG7o6tQzvft+MgYsmas
g2lVnzcsmxJxHBMlFLLKMMq+wCVx+K2OzKAXrDeret7ISryC6lim7HL3WpzGyfeiJO6gNC52N/zd
TWfetErSOpjiAAqOQxkUcdNchERosLQrHHSTEdjXa1zx/K1IIneDOwJTaisOEP9ar9vCl3Mbnjio
h0ddriapwmSSR0yUjMmkWoKsU4bzOHx036fl+rTSwkWR9/bYHPVVp7edIv9DvNF6URkhH+LE+bwd
i43lwQseZwoXgcmz3iWgW5rG8WgO9rSPb5wyncH14jCVR8q971/iWziZ4em70UY96NH+DAsw6xQt
mlLqAkQAUZ1SuOV2NNVDS9/v9ZZIwHtmd6D+3IcgFr2JokM4un5y0XG1FSHpJ6yKoAr6nB1GxqLI
yO9guQxZ9E8UgjYeijnlhRr6x+jIFW8x3vG7mEMiIrdjwYlYolbpMzzjgj9dghzd+AjnsmiAkRIU
566c8BEo341E1phKeslbXDczX//vvrHwTKpVSqd+OOMDIZjJYV+6dvUbCUa24jCsSJbcpCbF5nd/
g0uDtQcYS3EeDakY5TTXVy887LLWyPuWZQfpGDhKK0trmKkliEZJ6xvZbPjGohWLz/Lr+l+4W5jt
8SoUjDK1+Laul3vq8YiQsitMg9t5jXHpbgf8mpSneqiIbJuHBRKEdE6Iwpu/H4BjouJT9In9jT/z
xjx6JZOrRodaMQYB1HPa/k/sxSyqckxpi5fkgTBxuP7P6Zp3ljGIhIdnRB3EaX50mjX3S+ygUx1j
wJtt88dj0SZNajlCgJto7fMI3P0/f206rnEL6NODDK7DLARvmH6ZT5NxA7fGTgwUkH/d2kcdKDfy
NzWpYrex/hS3QHy1+GE+VCiLkq0O3PFeSRYxtW98ClOnTOqBamJaEGrnxO86xpuGyZizAejsifZ3
HPCfts7YqiGimrcnrff07+WwzCzeA/7BgTHKPjbXuAPMwilD2nsl0m3n2AViGFEkhKars4EA4yBR
zKrFnOHXE4ghnJbiAkscWgqfXmZDimPqbqHSeO+plXP41weWX3wRA+xOcvD/+DVMdZ6CCAIAtY6z
yXnqsOz1KInAqJqH7H5PCkeQ+9TquhbUUWGmJDIz/NCLC0vOsVX6ifeAokBiwEEZvpPm+F6sMSE2
LJOgzT7+nRXZPyKjWBYzcT3BKSuDU0ZSmDcIYAVc5YjHe8zSdcCfANwz+dnxqG0JkcBljvPSj6Ft
MWFy22ucm09lFh8ZctrWM7HL0OX/ip3r1sSAflhSrd5g2e2p2n7tmDZlJpOz+Kzune/0seh4Ay4D
PLFuVaIMjYCVXCNOjiK1PH00jd87QboJTa4zBV9VvuM6px4mTMk92fvI/HVmwoSrPPlH9YOdYD50
RF6Vy/rhQcHT0GPqPGD2lD3hYx8YnCTVJ9ieHE2c2JrlrcVmB5wf1M3wY/ZnEKtGO1xDjnM973Nt
k6g3IATygdbIX9FgAaENNMfwF9nSXqNHa1eQgo6oSludIHuemdptadddWDwtRk/JcTfZsFk3bQ78
Z9Q+hBJOXNaU2XY0Gt0YqzOpFGA3njRv3fIMvgyxXU23/jPCMZ9BU2vuZvvT2Gn68Y8abnrl4O6L
kIJJeMRjyeqpy6tWKvY1abhCXr3dCRkMQ8nqncUH6v6Xv+Vr9LxaI0+whndzx8Z1KnkeV+y5+enY
2e73shjh+iOAwyAwZymCDsCzMhrUV6yyLdMTkgAFaFffaDop5n7K2LqGWiBSUA2E3ubcIhJbXFnV
aAgy0ZcGd/y5AVMWM4mdQHnNxV7lyt3s1CKp4tXHziTQyxIEf/+h/SiOEUIaWnZTK/hR6WF9ARvP
Gcno7xWjpqMXPMVK1ue8KpVmK3uaXVGhg8HskEWcvUfI/EWc3R++FEHKLVN6bKdFSly+90XOzZe1
ghMN00R5SEFjl8f8furJ2ZtyOh8NIfVWzQAhrOAE4AwRH3dNajHQ2+v7MqYwq/8KReKbwANOqdnx
Ayy9MsiXPO14zZZKkvN+znmrYHw7Rb8y7zufWVyzy2CmyQdKBlRcBlbYKc4q/z2rjkAiRzcVvdfL
f7Tlujk0AUV4kl8CQ5Mwr2jn5whfUIuALTxnbo9IMi/cB3Mn1NP+65TJiMEwrfNUFJAOC3VdKy2X
cc6reU//pXUwwo93Jn5hnR6EISDPHEtlvJydS0Sb5TX/w3xNwr+qKCRDr7fRIFcgyAs/aRsHz7OB
NGmkWqcvu2X7BiJZQx5b6eE3JN8ccFQ0d+q0duyQ9EQ1e9ekDHBQypz7WHp4PVLRX4ukdPM++Uoq
h5WlugcaoD9p73fT22JFEa78hV4bBSr2NmVu9m07+lfCYxYmJEvziBaRpAlJVV3UIKF1CC1rz1cM
3WSMv+ttW77gBYkJ0HbtFefX/nmctv4e8335yf004SFm96snWVTlat8NvQ9Y1Cr3yfgKnyv6Cbpo
3S76CARTFm7rYBxnykBtB2bbuLiprdg6fWUY28hOJyojodbi6MIWLzlllBGW+eO3yutTAwQdmZVp
8q48wAchxHsoeihpRXfjEhIiawwdn6/Ubeu6mvrczzw5Yaxbz8k4xO9Abtcreyo2v8RqFoBe8RX7
KOpTtxeHQ3f31M2Jc6j80khq+U7zkURn1gBtsOx2bGZmu0b6bPXnR3KIRVQtBLObdi+h9RWBTVCW
kuWQKVShK8ZAOSsUgBgwbDPh0yMxe+uSOEHWqUo57WVgIA2Crtd5NYFnrP7L+CHx7oKl5plu3ykH
uqRZoTRsimKIqJ+bsaVzGZXOYSV32xpqI40435jBj6H+jQn/mKL3c4Ku06eik5xcubd56+idVpzH
3Y0WznWDYy+oLcdX8Az6y2K9HDzK2nzf272OJI+PVX9ddfxMoDmE0t64lvN5DMNMiOq/6bQ2fMB0
7cRbNZTC2QkPQdQIYOomdsjLd2NRNloHVU5WTeLhmx+M9NQYPg5gjHSSYMaO6y28gwugiJkS4t8Z
b7QfF+n0vR5+WgPG/6KmNyrFagSdFe0RM1VN/VeippoMt2rfRCzAjOW+dsMOLm6WK2gyGd6lDrZc
lP+fVDE5CM22HtPH38geVOl0nJH62pwVULaWP3AYTFfdpp21rFUXlqh1UTSNTzULbVSCCUs4yQBT
bNA77v1nvr5lyfbofyFGmr+fZRMqJ9JXTK4pjvMUxQJtnLyRK1UU2AfHW0IGwlIvlIngua89yiSZ
zo4iHJ8aHmiEKDLwqTftPLRYS31d2PZTgYf6sHL2/QQfDKkodDbhemRKWlV3un+wYS8ModNpa/pk
mSapMl0XQToEkjaFKhvL02UcwxzrcuxfwgKWqPCz0bXIZq+LX2eL26jZlAmN8k+ivsBhiumZZwNz
SAVN5SerEXjazC9dxDjkUn26gEzksql5H2WnTK/STUn2Aio1Tr6QdmbF2xHdzCgZqU7URUDPnXm4
IetLSOckosHAvt0jS2V0nAzthASoh0LofTJwFSXTTVggfQmTzW/idAsqF9Jn/lT5h9rXOsXqDTA3
sEwBLPvQfzUVrG/On4qzMaRcvIetUmsVHayugwG2w23sibzwIp3CFtUMm57Ll9FKOo8f5jR5YLHf
2bV6ngfSyWlJD7ZdR9Th5NPADrEUHWU6GNN5b2YD0aHIc0BlH+p5xquD95GYP6l2YS09xxHPGbeg
8FtRojDgW2rG90nQlPPGygpWnlMcx54448jgDVJIS1GArecMjcyNxCHd0isDjwAfFjvY+ihXZhRq
U+PosyMSfSDC41hR1J+PXMAXc9hae4Ns505okM6zQ8R46gwOMrMP9hvEhZqZxtoo838WoOAaBUHV
QlwokGAeIjG0mBf5lQwuNjT+WysLf0EhEg0zADj6dCvZYGzkbg0WnlIVh7Qjp7PdFmSVC9Gs1d7h
+ylDLG/SeLq6Cz3YJqhmXx5mvNYSlhQCqjya1w3aI51L9qHfF/IQ+8IW4PZkj07SjgLNF/jbkf7N
niI/5rRkXgmcnNOXT/bIyROU3ABVWgEavCWEDAkm7ZGKUJfg1hRxvbv+OmeD5jn2NHpM61GyhGzh
idteq6/tI2C6jIHuaqtNTRMzb/BpFUhvdbjBOiA1RpaKHMYeeevyT/S33vx82jnjlpEHq8bcXAuE
kEA8xUx19wXPq4cs15QauUjlcYBpRdag5Lfr4RnQyfGWnMZ75m/Sz3NL6oOPJFxQmCaVbhoz+ayy
ZW3IBcJh7f+AqaT5l1/qEtVUwlpFWAdyEBaS7qelIjG0WarCkgnh4UcAAgUEFcPuLCB6cGOk9XNZ
apPv3J9reVOE2CHJj8KlXEem/ujoKPmO1E/nCP6ue2gQBtv+LdiulvIAEBrsA9avi2BRsnN8rTvz
4Qyy6/jQ9IcpqLwY2gjUbtCTMLRkaYLF/F3qYYa1hIvE8lNp+DU77jFS0H1BY3jYtNIJUQQw+j4P
0lNAvWTLOlsTPTIh0A5M2wG/t2gyL5NTN1yijMFpoUxeiR9MxbxbZ9g1epmj/3nGqM+9wlFQ0ixU
TtqYXBCfNJYxUFbXVLFaXauJ93DTCmJAgxv/MwuL62AqLakQag761Cz8bcaPxbg19Fz5h2BMg2vr
U142v3VE5Rp0maCPZl6+rDD9QZmgzVk8+5JXgHO/jCYkATBwIkbEbd83xEbOVZgs/4ZYRiwEFFVO
Z0kwSfY19qhLjzzUzbP2YWv2IeN1kSrBVs6l9MscUvfi6pH8dKfVg1Hhcvpw3UyLVOWv32BDAwij
BVoP2k/5RvbnHri9BEizhbvf64ycQZKlFCWru/l+O1FDilKkRQyv0ttB6Zsx1NtSYwSpc+nDIUkl
akdy39dKTjHNrNUbgvoQ6GJO7sLlnkgp10gMPfSVNfPjTW9eySXvFTwK69Ic3NZUVvqjZR6dL7/j
DJpvz4VTUz4i84/CGmV/EgX4H1YJnEbr0nfvpRT0rmH9grMd8SI7w4teqKz/Ok5C1kmiaTUXrhfK
d/RN4sMgyho4Fxv5jq+tMWGiKHNFYkzoHZAM3nSOEemSW6UT9D5LU5/u+nmxKuT1LdcK3di8bh8J
u6xHZysD5f/tecU1KFBsb6/BsUjqXbz7PpN9gyF8IPWOaozHyZHJ/dAHr+BleUpjCQMtTCxRTk0O
kX2s8UnQxK9tG9KiQh1Sadw0/Rgn11VYfIvR5tOtRVDtKTui7Do9UBZ4C+0jVgn1Ur88aAMgSFqm
2qYwfYT+yRwPUlwCZLNIgCHBiQkVtHL0hLKo+tVK0dSzIicG+h7plqeeipzLqLOC/MJDMRDBtl0Q
EO64IDEw92c8MXqHNXgYET84TR8jTpDg7yGbzl6mhhHrmy90zVdVckqQr++OeJoZsDI2tY9OzOYS
Z3RQSJBoKbWv5n5EH8eHOdNERx2tIqzjCD3OCOPWPQLOahlv1+URT/FOcYc5cSoZMzQa2KqkKrgr
K9/MELJmr/iwt/4BeGD3GuXudTNmhqfd1kiYL0a98jIaf5mpN2HGaC8vWVC/hWkfoVtD8Rkf/vUG
HVQK/+KdbVTbRXP9+s8K32vUCyscAC7q8a6orWvH7ZO7VdGO0r11mJrNmbjAJD/Z+szGHYQpxoeX
Vc68U1U9ivbD1P37lg+SDDuF/Cg6xrAcPsBem1SCl87ZYWJf6P8gHSSVH0KhJ+JK74/tdfzboBhW
g3KWMROebmxVU6ahCAXZdWxq6D2ZpTDItrIdfRwRdjL2HFANEzsQYFJqMI5f2jwk74qICVmXlyrH
P+1GsUy5Ln8+AYKw7RJ7X8upoblzck3zwI4a6yX19OoFypKk8xFtpbpVl4C9i8gWYa3pp8+V4drq
19ZA3y9WeMAe2/V/2OtVBhRN9sGECsK/WFen25wVfRhJZK9A1mmTF2mEh36PcDQq8a44bNlAtT6q
KMp2GJO2YmZortqG4aHBEdbr8UYfI9C3d2xvh2WuqxImcKQaSJMyML47v5tfwaLlSLrpC9Tc0txm
Pq3Co7U9PJiX/j1HR1RgNCB/k5DnY/4hmPQU2c9wS1CffmbTrvJhMkT1rvcbTaII2gEZ/WBDAxIH
A/8DRoPdPwkSg4R2TSIZDTvau1HaR+Us2fqH9AHKE2nK+tMmTEU5eSsvOUL0TFb8lBXx37BwktLm
LVqAj+RUKFbpnueuv2rtEm2yB/3fabAXl9mxFrZvWJSknEkplXuJkr2HxobpRjk9dJh4NFkZu3LZ
+g+G7p6IQWvesRRvXPR9yVE6BXh+lDqzF/vkAL1yWNlv4S0QXWkZilXF5127U+52O7wlnL5OghNb
CMxj1+7IIMjEMdkvKnccaqspd2jcro3VVXFAvaNoyfLe5Op5aMKtLHPu/yr6IGLdv10b/RRRh59s
hALuZKIJoi3Dxjis7oaCu/glVsT90gAEEvk2E7fqJwckjkpRZ7YJk8z6EoGuEyt2BF5tZw70SDtP
gCQs0Mbw3x3YuYlCjEiS9B09nci5o2gpMUN4mCDKJ3Dt9wpZMyaZAP2H9RcOxczjFnZEY0OBgg1k
qaPe1FKFtNJ6qi9VBTto+L1Mr5OayKNG7fB63Ku/oqyEk9o387QgZN8VHoM4d6QSoLE+YEriPuDd
5c6S4sUxDbewvpdjp7atGe5Z7q2TxMoAGzdJdrIjNB1JqhlhxCK12HskHC/qYMPgrOOm6xmhC/2f
f2xtUMkdkA8nBHTurhwe0WL7tU6r16K785PI/DzsgkoXm5axjQgqTmKkmvVUh/IBS0Rs0FC8dX+5
pIaQRfVGnIBBkt6ghLrWjoX9vACwbM/iXxk9lKMzqR09sC8ChIwotAKYfRz7EPYYxO4BDfOFJ7+X
dXL+5pCPWM46z5L3gNi+ArMiJvR1bqL6FlI4lOYhnCo3EFcCoosMSRcEubqR5ex7MdYRbgwGyiFi
Imu3VSaqwTGkdlQEpViG+ok1GzjtVIEFBScaZHzGieXgi7d4YyVKPICXPoyDFiCLuDaOQD4sTchz
XdUD//xbPGnvwSfuYxGtNO1ifVBxVUIn27kUQuENT7tepW3mrQZa3PDQGeYSSZPv9FSs5To35Vsp
hTRA29AcW130SmFJBL074i7n3qRfZjt1w6w0uPc3VwQtrkA18hyfqsjwS9acmvLsMupL2zneUk9F
HUBKJQ9o5OfxOdwf1lWVGSBXH4yrhTSSQRjvoqzo2jTWPfQwQRCvFcFW+fpIYSGI6/Qd8E7pf3TU
cwNVwk2FoaJi3CB9l7RM7HDNwz6FxeogElHo2AzQuGFPXQMj0XzctNfwRrmyhjMFhtSWPiHlFVap
a+r5mngxchtlcilOc8WJgBmS9VeOl7V1FvOyxjQu0L1VZYTb3+w8l/lbthtrzUbkA3v+6ejU5Gx7
E/e79lRed4PP9xX+5NF8bGtpNOJYN9pZsq99sqTFMz96ex/duQvZQEe9XyD0+Gmi9/8TxEYFsZf5
140KIfNnyr+QgC/NWHDds1DOVUqkN02cHEaDgY7GOdZADJNSQ0v2/nxz2VuXkOVj56XoiwbMtCzG
yLOphaSA+JvrPvN5ikJuOFmCTS00CaALvbU0jXV3PQat5w+5nv5Ya+rgj7qHPv4C1YdDjA7OcHEA
AT4RAxANdvVZwssx+fxj9UEb4+qMTzwvNIVjDEbkQteAoDGo6a1qEtE+0mT/poSraGnqvI9wKbWI
yCM/UXOVboVshFXWfhvhHtK0xJzsvoO73HR9NUQVigjOeETF+gXuzmRKSJdnMCkyqECoNJEoWnzz
4/7zvRZW036DwmOQAxsIz3E6suoJcIPYy8bHRl2KJM+Oi9Hkt3xvz9q/GSKTGjC0blJStQHVCN09
I6U2g2Tfabfxmy6l0tHYI+g5Wn2RQnyRluQosSnHMmcxOJXQrT5wRA4TeVyFRZKx2QGt9hniQIOm
CqAHUchTASxtZrkOQUAjjtY/IyjDzzsj5AI1N9cPFhPRiKmm3ncKoK3VzyizoOT6MozcE+UNM8bY
710PSy6ZtESAsMgNnVybVDdYRSL2ImvOwGnHPfJAwaiJNVN9ddPgQ52h8hY9nZskuNg5NE8c9Xjb
1K3QU2zYHmyB4YBZnJcM+F6t19C0x/Mx25plG3iYHZOgCAGpJJzCzrtjl/PE9OnujVGebRowOapj
hB0sieMb2hNGvLK8m/w16SlPGJbHd0Ag+Z30eJwS4hg4lHPVCL4zcIdlPe/GtFauhFuQvLw5c8WU
dA8n/i6kJ2Wgigx7Ztt8macCw6YqBN2H3sG5d6OuHN9jQzSvMXIUyoKSgFpOMk1XfT5paimfPlc1
fnzMZ+sjFybCIAxBcZNWUJpo5ldJ8+q+Cu2DYCwkg/JUbZBtAyc6lJlAw0wiofZJQd/1uaOiPL9c
UsJVwLMQho669Mh+d4YU0QvNf9rQjZyPO8A3D2szbi7JkIZEl00pD4crVw4gYV/P0v9zzKte/Ixm
5mzmvLGNh2boA5wFntylMAgvcdhcKKiM/izL9SQZabrJGZl3m6vWazNjYRaOgIL/PgqoGgUXKB5U
fqGymGOBrfTAX9TOFOwjZweaAt9LuZaMFfwI33vYNUkYA+XNwPM9lV08ThDnI6t7h+OP7K42J5Kh
qTUez4r40cEjNfQgcP4SIiqrMd/qu0a6lvKuGEVEefoBJUCIYsDc8p7j2yg8qNHdiBgw1Ndok5Ll
wuPVL0QwiVJir63D8pW34CXifpHWshdW1WmMnUSeWWyqxXu2bEtC2PL2yH5bZtxmZrJn9873e8gB
jU/VFFK7onDdK589K5R49JIl8itW4qwXQSwWvLbxPLHONQ4HuJFLjslfWvVJRq2qt4BSSXO+TjEA
UXyrPx4nQ3fc8j9LPv2d6TFqLCXaw42KdicdOfruKdbq++XYTdGCgarBquQOUZqsxTkRUv657SBr
UWbfswOe9aQt3ylymlqzlIp5KhykjzU6uZ1mG3zTASBI9zD+08/iGm0SUPTWDhN4tqnwwTp4dKSh
xe1E+v2wh0Q8JfTvof0HeyjgAnj3jlBYu8oiTQVVayg4cQU8iW0BtneLowAhWhlh/QPg+WvzFnUs
U43WVFrMO7q8GRn+nknyfFDTDncwAP0G1/o8ERLbzMMDoKzNTEoTc6MwFLXKMKZy12AVMPcoPmc0
L3FmNkc3Ln8ruYv7PSf9HborPBpz7bGN8BjEVk4JWO9Q7QNFT1NUrYj9sLctjaCA1sPAZci20U43
INx2A2dZqQCdoYmYeDfW19RVv7dGxppiLafk5YE61/WlioqWwqN9s7evBCyT28BTD7Mrid2Gqe/6
LGwDiKrYYyD9hJ2HFcJau3mW/z8dKHXd4dwr3jZY+KvSY9tF3Bv3qDoi9Q3TfBnihkiE8keEC98G
retQ/LwU47fHG47NJf41NjqQUJTwCRwFnKzxsXCRTEFV/dJvSJ6+7YEzPpPxyv1BBmY0dVY6AucC
aa1aFRopqaRpPL8ELSx2YC0OePO4q8hmW5zu2ssdwKxU1yyqIO7AT0eaWtSoD21/5/xitwspA1LQ
GANQXkXZdHdqHZOuKq+/3Cuq5dTL6p+Ns4Bk45EIoM6Mu70ry3gN+EUFLne6P+GnCkxRT1z6znDU
IWKgFCHAiNQYyg8z0mBYNEri6Jjnm7vUeZEPVY4bnj4a3xRg7KQx1a8Rprg1Hkui2n8+sQnzPUgA
O39F++3uxkmWiQuYw9n5Ps7fF2lXuvad9sV9i3JmAAjHj9LU0p2j7BBolw7KxHNhzeRNMApn1kGK
wInyGn7RInNWFX78nvNx/Dubfb6css0lpd7xsoHv04dWKSL9U7Llh5PmCGhEoilbSvQYE6Cr3ACj
Zc3pUAxZ+wzxNg1PuILk3UHkxkM9Vk9JZ7CLxG7rfwg/HOyIBCN9dQ/3MaotPQmXVRq0O4VgURZ4
jO8wzSRIugsykweTRmBhk5MBtJVs5E26LSalF4DWMBegfYeZhjzx9MvBR5sp+yxWCI20CEF6S1D0
Ybt8MDlfT1+a0z+wwRYz1sWjutXIp5Ng4axHewXVqeD+nY85HDevtXnROlH+Vyv11eSh+c/5/Sob
evuaKvJYml6/Vxpt+64FLg20RwpDN0UiTDnlT8IO0gOljBfHLvJARUwlvIQq9wnBj5GrkXWfPz+6
d+gAc677SMpTtYpmla9oj3jumNNnIiZVkgAGGnMAsvcSx7JooZduEOih8LB5L+JMfEll6KcUx0GL
l1w5P8FWlLA3dUA2R6ybWqxGSxO/xTUuJiz7tno8PWWbJdvDYbs6tHOwKTFUoiZsuNU7sXoPLS8E
Q6BCJIId0ceiwqbkzPJZeATmxpz/OVu48YyZQV2tWcPNcT421h4oTRAdjHEh26kiKGNTY9UAPqI5
pcrwNa5/js7aTKtkvny4VBWkusvnZiqpWzMurQZM1ZNND8UKSvUhIu9yTF3wFRiJqu2VStcptDTf
ULTq39gWd1zwz7dQxn9xybmQZ4RnhnFz2lb9r0um7EEIzdauoGjjXvFwIMevDp6TB52djg/AbT7D
9MF05OlKJ5QiBCZ4UQE+gfcNI6nJjxeBTAlR0wBb8uFpeCNDATogCBE3Agi24p+gGrsegTW3djVR
ryYhuKA4EezMFxKpFr9afKzhm33Yfx7tE1TeLP7GjoJ6evikNKppJPm/LctwWe74Te4n/nlHkicV
iXiVCCQ82MJhqSSR197zpvzL3nF3ji3dhaJI3QvqB38T+J6ZsUp4oRBgpKxoYP3xhIEmLQKC7GUb
Pn7h/9swOOXnOtThmSikHRV2dDkZPQJ3+e5fW07IFjtZ/LY9TAYPn8cautI0PM4QJL6F4iUSnwDL
fSF9bQLHDRQC+eJQL7+/uDkJG+h3uKNJJfXrGiapoPkca6xu0kO9/52i4XGaFlpNQS+YghjerojG
BzaU0RFiRkC5VRz2rQwaCsFoI+dtENKw6Fwvp0TUOJ3taFzy38kFm61/CZmDYHZ9OeyMGdcvanIN
OKhzWHyRHI/kf66jIHE2p61h7s7/BEMq1z8puWev/j05cogKspwx/WHP631hT3WugiSvN7zDNmt4
MuTw1MFpDZhyWJD+sRuAjVHIbIsYIYC7Jc/sGF0QeWwGnCVL87ZfxqUHI3fXadJSGl/mRvDSzPlh
5bC+PnVkKFFAXlVJOlEvulI+O/Wf3rz7FgCNcFCymGJgj1NgsecZZGLpKgxkwornwE/nT7XGNJjg
vJCrspwZI/TDiqMiINTtTnx4loG3MH2dZc60SA8cLDN9pftBhV9+DO0a2NdnnkIKmjbNJrD+XwEh
CsPl3tFqgGlMBDd2INcSNefKFtCFzbsCv4iIWjiMFtnnJlGLOSAkA4iThnT9ffeF53e9AzvSntD7
hYzAXTuTGv0ZinMVNs3cuCxPKi4LQsQDc9JmcozisGnMSCVcJGTtq1m25j59ReQdr8DEe7CDjnLb
xyOK8cAWDpwbhpi1THu+nc4/Ri+KObQeZlfxho0j4AWGqJ7RBOgOyfmTs9lcjUTX2H//TTLYl5BE
r/35Vj8PASf6SIiJtq3Ga7VXRAbHLW0e8KDa97LD0KNSpSAOUJ2ENtI8HASkEwgTcYoUd/21542p
q3/V8m0EbdPToiJfLHgrFaGAhk0ODqRrxwo/KNRmz9cA0tneEY1mjoSqQYDCgT7XHS/GSE2qSr01
HZC9b6ZLtBvBdcIg9dTLyEBdJAEQdXk5IQwYpKbE9fZI+FNwr4rTDX5KCYR/1HRqgnZ7tDklhSXP
j0QFZV3et81TDlmqOzCA11Es6JiECGrpJMAUwIgoDZxsZo4WoR59DfkfeASlyYUhYI8IyaX2Pl/S
9DyFeRJ8FVC0sf0pllxOcHvew0jqb3psMX0r23Y+ZtGTEdnyFgThjqgWIjcd6iWHyzTIJqRH4GwK
3rvNVL3gE45wCPTAP5RqnKqAnTcWBSdcDsggJYCmMeB5tMj7kUfzaBeuV/Lwvmr8mYEnvrv4jP64
cEkWggwa3ebYmlQnU464bLFI9PQU3LNd/WTYUscS8i+2+a94avSYEdFPga9vI9ofZbUI2wCUPuUM
mqUfUb44tPyX+37tDTAHF7r1INB8nW9pPEoCvuFfwwJv5fP+T4e9yl1+m0xyCCxcDYJ/SX0caX3G
VaZEd0tu1skY6CyS3LjXA7DXc15Yl35o7x3D+DbshNdN44BABqxKjIOlduQkWu/BrU7B60Bvh8pb
UY40+aT3rGpkxZVhwXykhOV3Wabhr6ocXS3Xcv8FAMH9WzfzlLN43t2idtAhtCdM5F/91bdHhRV5
bg26WrdZsLC7bZ53e7w+D9HtCLYZa1rKDZVlinlTStaVo8arloOi655DLS4rVU49pv8f1Vzvyi++
RQzHHYXifHms3uWIGGylv8GFIfvqSdgzT7A6BolaG6t/SqUiHhnB2sKdDs537woOxBMEiYR9qvpj
/vKFgt6/jsO/T3dWgybSwr63fVqH9YuUr8VpeMx3zVq6FXvwKN7LOrxk/mWqtBAYpQmHHw6LbAvF
V9SWmBY/CESvyKRV8ZYIfeQE8onevsppxe4XTnSWQLuXBY5Wkmuj39G40sU/65kXsdAnO7LmzF4T
e/5R71UcU2Mvc4/+Hn8+sxUVI6z3F33c6XGalkkt8LwuA6xEZORvGg1mT6+/6qb1HzVyuba6NH6h
5pJQQTD7hiR2xIibaPFWFOH/I1y9+AROCbXa/t7/h2GEM+nvbxGnU8FeHYkYTHjPQU9uFFbJ7coa
tpV/99Ug7eGlr7gWAZnr/n5kEc1/cv1u5Xp32PSBR+cYuVeljKmVHIgZ9WcJ0QyAUTbgvxYeK28T
G4gDrMSTtClw9bnFMqfmFs4ajDraEkHwH+4jC+R9T+tsKh/N9TONa6y4Dz+/LaFzAbVrWN+hsMnx
aT4ZmAt6LrJKm824dSeZxybvHTl6F/9fUhRnUvqhkxzTPGRW3Qj36UBvBf8A3LaeRcdvxdkfDOQA
+o/uBGlr8l50fzpjDWrFbqDaO+QRY2T9U+qZFO41QTT7R7d+cLCrYp1Er/w10wFMnJeBigw0e4EA
D8n87nRFQFzyI28oDJKHO5lgorDzMITgEBtaqTHEPAquh5nfrkPCjkNdVWn+PTi3ewP+6tmt597j
EnJKniU6TiibVUYv7ehPAFYtgHc/AXZdvQ968oMSBq6Pb8bf62YQ5AJsRNB2YWJiQRxPop8JsHjw
WXVmZYbWogrXsleBgTf04aGKwRvN1PLpPlQ+K3k6XUTB0QrQbgE93Yldzb5kkOnq4HJvfclYP2bC
4XTb2dUA2TZsFuV3DezZEB9jNA3X2Mtsr4vMMWGGKXcTAAMwJXU8ZsYNTi6uZZehZeKNRFXPTser
we8gXVhcn12VMphdxYAE6xskc7ExQbxOFaCu6RbZH2v4W/SA7NdgyQEYvJj5IPaTQpWOGSFftZ0Q
KW9q7Qq4Nn8KnxuwCU4mSAXfwA58tfYckkoCZUzF5KyyPxd+7c/ZDHu5FeqOSvU8uBSTvz3BKOxC
GfYxbR6hxAmnmJCazYzEcULOFkiqHRU9M/eMMBgVoc5WcT5GGYA2837wadzVPSJzR0niuM/IV8O+
jxkN8nCkzT8lJuFtM9STtZePphhD68/hsGNj9OPfjysmVIEMOIhwbg4oLM7w//KvpZHd6vPbgDkq
349TQkv9YYv61O4U8jOTZg3KE9AOfvdLCe0/zL2R42iCEEbp6i3so6BW1c/B1tzdH5u+ar2LEWsL
cqCnyPdTd7HDUi70JdCl7COxCqdw6l0+gryIDHnScvBd6KKh54CNtzYAS/BWUuNfCbvm6gMu2J4d
4SmxA8lgnZfwononxc7PMzo49GDMV/1sBffIHxHDOAPNg4msrqnTu1t4dH29YpXlopRGUoxeoEpi
BFRm071ICR6lCq30lQcnwuAlG4FcC6htTErI+rnhX6mb6S7xoMX0v+WRnWJc8Ccd8MJyufYPUIWx
AsCRGXPzhSMfit5sf6S11J69MH2G8XG63vw+knjPD+qlhoUkrz2aOVWnWMukJLSvAHZWjETzOtYq
bSnLLg1apuQlMu1hhH5rD91PZ22lIffjaC/z5lEE9jKKbww+rbWN+GwheirL67G/nABkt5bUq0X9
zI3HJkCB6nEcEJmZSaSDARE2JX/Vdq92HyZ+XhieBcM4ZZeStWegCRXjaflNnGFnjikuRGXBYKeo
o07QXjU5NkL1ZW7KeW8BBGfSqAoDFSpJlDDfaWDgNd7tk4+cQqMpE3Bi9oy0YJo+tsrEfF71oDPk
ZXPVVoLiZ6lo1hW0f2eOqtMaLNUw95lR9cysd7LwJcTyRScwJg9DTF1afxX4GlJy3+U77OZrVKJB
IvDKN//+i8vGtI3UMjOdb9JIGkN/RWNfCmJSeVMnxo/CoIwXkW3eLa+pfoJmZkAqRAkaG4PRsur+
phe0q64xAJ4mwuBoFcCJ06E9YLEaJCjW/DRR0ylS3h3iY5RysQUie8kPOcTyrsI16Xl0vuLcR1Dc
36DfJ6K4W3kD7Lojv2nnp8Nxg3CmNjOMWW1Mm++9L/IndizmaONcDAJ/AsBWbnuFCyMqx0u44KeO
NaKZu0i9BKWwHklwYehd6YgnSrqzhkCegCT3Bw5YO5draUZkbE74ubPRBJ2MHK29FO5UFfylSflb
4HEPPHMLlRTLPqEfBQ4i6rdl5HaulLfAFV6hgt3gLo7VYNMvZIn7ObUaLn0+4fSxUPPR14r2w9P2
wvGHQXV44jU5h1DaEU6/nDZwwWQCHxKNjZe7lZlOVT1zecTFTlgJkznMsauNK6zxvOwWIwnp3Arx
lhdp1EKlBNRCygAcGd7OqvViMqtzRAig8r8NsbrpGkTm11audelEN0sPgnFbNUmBtIA08P8K1Jym
CJW1wVDEtdbSfLC/Eplm+D0ZkEb2ItT0fRA4jIPGSRrSQwHe8qYj6FtgQ1MAvvrYIkuCSUnytewS
5VPNSNL/LK6Xvy5AVnLoYG2w7fOzCwsTBy/ztjylxdodXne/MMtvbwNlN3shmPJTvDVsLlVECkVO
qBl6EayGqGaMj6l7rLzaEdndQQhdZdObWQQIFwsXpBa0w2Si1UhtnFh5Yygj3ZdwpH3q5pXr+g6t
zekLcQMiKuN6NNF0PTa6x2PWbRj13qoapUJuly88olwt4+0vNEXvIeEcP/14V6YSA5vB0Lmq4RBy
XJZB/D6rFpo3qB0rXS1Hr1/QIOhwlAb/+zsdc/WB+bUHOBo+P7MnedMFhwVCGLPu/vSVDJO8TrG5
6/iOPPzAIqQZQJleN7hwd7nXWD6U1+g/WZ3GlapaIox01LaaDB3XQ4mOymjmJoyOEqxxfoCyDvsg
uEcAbDk7Ihub+JjHXyQV6b1UVqvEVYcenvo4h9MZQBbEbmh6HrHHvidqOO9o18nRMz5oxkdtVu81
fD41OGJl6hmpWXjN8bd6itQVvpTsdgYW4xilNGRHjI6zt2Dl3NGQyBYbRAy5xb8tvzZS7poEeS1Y
A4kL59aa4zyA3XWVYbX43sVSM5hsPc6/jexcvK4TVQhPVtkFgtjaGVNW0Dg8fJYUvF1dRHBmFewM
NpDjjGpDutXKpNt5pQBW9OKQPMbrcLaXu4K7h4KS9gVLGWZJNK23tala1qv9tMA6MsgVfVTpIMHs
9D3lR4EDeVcD5bb5ZagCKuMFalJ/EEjQaITq5oQfBKiMXge8YDZv0jrcMPIwre074NcW+nuQAwY2
dVD4cvg3IFqxBgUsCEaT5NaJ2k45zVik5d4uaaHY3VthCLtOgIP1cV9zSXWl7uJ2pmrCxFV0KwqG
qLCAAcEDyPQ+A7hJ1/42w/WYYEhNA8FULKzwp9n4OyD1XlS3MpuBBNDNMVAXA9IHh7BgPUo6FWgF
t8NYwk7H39OfxXqJMetw/lBnrSNTMRSDQknJk5ikx03039OIXdi5iynKzOXohN9aFq1lLqDJu1Nw
vh2YmuaEehZt0P0gSQki3GIj1AvrwS0VpdBpjGLtCT1JWNaSI0mqTGqb/JfmA3dPcW7NLmIvoPow
UCnTRZ9Sn6Sj5rXZEOvmvR0Sfj5J6U6njChGrCXa23UCIDDuAy7bChkluQF3elKv38VfWwU4mez1
jD8qr7xfgfEy+VAq6dPzZ793kEiXCh5Cvnqda61rP6jw/LZGyZrTCkuKiDp6gUU1NGiAuvw7CPnj
yfeX1rfOG3p4IFFwrhvbv1+d8YXlh8UPjDLJe2HOkj95CFN9uMrz51Z0Yq4mzrptLhwgXOUARDu5
Pk8nG0NVYJTxv/wRHrwVqXBrjSfLVxLJ8OOPBJRcj0kf2oBz+UTLv53BKOL2wfzUJetrIbgr7WRS
TjB7W/Oc7358BOG07vZTatYjSt/oCDySSsZBrlnFnaAloojSC+y/9DH1NknuVdAZewAWtbb3FPy9
od1sDjoTEYGgeMVX4HL3SRMhO7wZbTSiHFDzqBOj6K65Y/Uh9K4zfegfEMa4FKDQ1YNgpVMZK3yA
aaMnRuQiLwmoRR7eW1x+WTtHbdS6Jqy07G07wmY71WXIRYyMpq1/KlQH2gsSUpCotwwJH00s18dT
AUGlcFjYA9wLdqxnv7Z/1NoV+yRXhOiSBp377/AWPNnwSMngaRKVAcFCQ1YXbFyFWn6CIXFcS71f
HPsFvRPjt5RutW36DrDvKtZ5lZ7cWJc5O85TZE1/m7zRCSq0y7dkdgRORPcl1MHlEjP7vAxcjXUg
g8aHAIMPnMuloqq+5q6qrbqfjI8ZgOJs46wwciibxpq1qh160omngXLml2TGYuc/TXR8fXNs0A79
fsVhKDMHj9koYiAD/+chuWMr8mr73lP0xolSCQWZcVGNumHsvAbyWmo+u22TzOypOP7oxUYJt8Wf
DERhq5tk7R8VS/dt63ay1c84u8QerHZ35hdjsAats89Aiyx8km1N4dIfytiPzeBdafZrZscLUVbC
vWy66v/jG+QVdyFlQNUekMGC7Eoci+W4ZbnWeUK8uay6DPRVRaw2O2xK3zm9Mt5MlmOxNWrPCcE0
Txl2oXp/NMPDzmFkMNqAHSY4aqucpBuCBgmRJkq1kb1a7PUbgrllQ8Hn0Ht0FZz6u3NpELl3cQAp
AEBZ3ggZk+a8o2ykidIUyBdXY4FWqkSlMOWYpAXvdutaJlDZzjE4r37dMeJZFfqFcrR/dWUo8Fzx
uporTY83SphHQChN1nSIcMZYVjrzjcwxky1IeV95tbBoCf4hhZBFyS28DtGLWJTEmixRWx9xeQf7
ErFjhHrkGD0QUXiCsblLDVbWvKX+0R/fSNuAV0TtYXU6y6nNVZ4YEEHUBTc5K1f7rcQfsAni39h6
B188i4caFymWI6C8RE4CDXkFJ50FXtb2n9LyPcl0JUMEx7Z18sS6ttRmigdsFnrvz5JWHSDeP/oO
axu1OP+Y5ObOdMoBWatAyfVLWfb5oqG0RPVxcEQ8lzgVqQGSGBvLEy019BgTQepYkgnGeZRtLfGi
CqZdILh2QYzBu1cphszg/pAEaCINHwsAz1F/5x5MlEhaomXN9HTyp6xmPx7kbwegaZ2JicdoQucj
FwbpxET+1aEOOoKOkdSRRlbE22XL4hsvzwSJVDAkyAwhKt7vF5t5jjjhKnYEMZh5yqKxRdop9A0z
ONekS6cBNJwygxikPoQguo7hF7rLDX1jdOmL+POIIxsTT/oQqnRjPlEkHIX7bU47R49zcqyOeqPn
uSfdFaKbTLVhaGeGDZhub3ucCqvp8xih+j9PwBjbeUClsKBukavXH3Z+ucwRo1WFajYbRQpCF5kC
ZHy9qCeId7U11K7b4TIsVAjfOofTdykUoN/3NAn9AwHB1679FHbfKlcKP2GBia/bPTdb6/DXZm7H
5XF5Em9dUo3QNEPbXrTkaRVARkkowB3S+geNlPSpu7jwn1GMtdjqHO+VYj4wXwdt1EJ4F/Xk0mPx
idDrMq72qurCZzA+Kb3AnkzV3ph7OUkpt6IOdp+0wyLrHfse0qyAybIx9+LvGRraDHxdV/Ir2SPb
Erbzd7urbacqnrrpcPRYlhb8dx1IU0uBRETnn1X0//6ByUQxU49VmN5Dv3Cob3odpgMLvs/02bNi
aCBBQsGt96O4jjmUCb8aL1gn218NSBsh4yDWQTpPMaMz9fKTt+inZvvK25fis9VMBN1iAqlJCZdM
94Q5W8mm7Ks25j+XRuZXNw+NdvTHyhwo6bCsnqPd7zcphC8EWkMV+boFfe4na+/KorV/hwZ6FLtm
cmp419N0b7c3fi51BPEG0Z5ZeLdq2wx2qPi/dWtBY9IGW/smygPKLjND4cXwt4ycCi+/UyViAeu6
t3A9nrzKYmnvPTCB6dsYnm27Cj704VSu7mFTUpm6+8oFWz1nIo6Jss8rZd1N7UYj+B6vH/DdbMCh
JNS5ZOxOP31NyILKDYK6+PumgGASwA0l6o8fZWewiKX33mQVHdWAuK2B1NCou0UiGPRROt+2aGiJ
aTjHSAkv11OlCbPjsLvjEaUIiqJn7LxmxUEKAdreoCxhzfqDVoew23U1aEfpHLAMPGGq+zcDhemP
t3DUbCYXjxacyox+blXbVb6cqeAs9iu/3TzOwLFyq366wMQYUPh9UFjeGRVIUctx51Ua7L2Qzuq4
Sui1MDZA90fJfIuRdIp0duU2I+ztvvBGUKsz8iC79kfIOZo8jNryTRK+tZPfMzUu+zkeVtvoEfR3
VKY58E5Ssz97JY9tW1DBIe2U4H4jpK6eJQOAQ2xel6Rxj6x7LHNE9FtVM7we4flvCklDi0N9qHo1
Gqri6AuFLAexFMG7FxHuV0Q0XMU2CMq+DgapKevZCQpTb7XaF/3m8Ubm3HmGjeLINGfVYo9o5xFQ
dtdlQ5fFIfmmdWuGS6kYoFQ3JdkJ+Bd6sFbDryDblphwEp7nUunZDir4APepNbmxm0fv/Tu2TEsv
Dif3BsquEdoWiFu2DEM4yMjqH2lNwYWGClruTCGYnNKFXmQjoQSXBaB6yY5Uj3+BnlyQZAUtNweT
jLjJ84klDlv0W/+rs0ExNbyJSLIXuzL0tTWBFSWztEI9ocVQeGQOK7JnuOxSTlcj72Qj5tZiETYO
jMg7wksUISNdPDRGen7PeZV08QYFLvpmYc1+qR2MfdOqtrNbOoMHxeVrAS6cO1JZq5pr0uj8f8pO
lJ9qI+bAA4qd2DS90iJqS01Rz0YRkMYfmRI9C5RoLyzz+Wheymag7XUTo9poQCzMf1XDan2dyrok
XYDC/z18RMKhRDcWp+NJvveRSNL/x5pJliPVRc5cYTKnTYMsP8VZ0xMbyu2GAo00sRxP9r7RJyTd
bIi0ieD5I/826jsY0a7K3OQCasH69h8X84SAYt9Ebo7WOyOE8USc5iU0uvCUerlvrBqLfjAUDaUD
WNW03D8JX7UV0hZzfs65ZWyBeCAH16NcHLe+djFlTvY6n1eR4YfT4TwDRfSx6UnLiAg0QfwvV2eb
mO1ny7rGflAC9rtZZhpN2zkBQ2gvBl70ZwXTLm0UglHgosa2SPAp2dtLGeuZrFS6T22yzHxt/8B8
zQbw85VCQYprLCu788bP3F4N+JRvwA9ZCxvVvwTBnXAfPgyGaXpIVH2pSDirk2lBM/EwhpJnxJU7
yaQ6qida1Cv1xv1DSP/JAOtovm40zmIb09Nt044IpsIUUlJ/v/WnHipX6Y0FxqeBuoNFnruosO8K
IxqRLdyPIF+oFeoEi+ihBESNlURy6Jlt6hjdCO6jBzlxk6gKpaYKneVMMYHKGrdD29Y7868Y9OXg
+stbvxsu+hMfRRVFFcsXtzcfU6BQ82v7p3ysp0b4JLrkFLQnF8p45kqaOZLqB1hJGLRZ864OnaUQ
wzocEZNL8bOGn5BtN7gbpBHw6aXV0lIF9vvqUdzebFDizrK0xCv5Ek1l45SEGsSMosEcWFigKPe1
RhFXQn1X6Zfa68KDQdMedCZc4rHVG7Q2dpADD+7/v4C0tgc9Srjt56uad8VUIlz551PS4yXWxMAP
GmWKOEq2ESkBFphWla+7n6Aw/EQukG6Rnjj9VNtIssprYe6x5R8e8WVmKowHtnQMAiJhT7XqQO6Z
q4j41nAoHlZAZ9zuDE7WSw/14z59Mv6iRqAul2V/TBz7TpIkb2T9Mst1OCqC/kBvz9l6wzZtyt6L
7yYTKLyUj1sijKqAZU3ASeKcEZ6bcCLBzm3fOng0S7tj2z0DnjEKibyQHJMkqyFCCw3EHq0cQcoG
Dpy0kEWp4Ya/xD1m1tx/xceA0Gnm//PufTxOwNS8PiEZbCmM1ftSPoaj8o5TcR4v1JX2TKjcJ644
no0Xzjwd7eD8CyihnDBXfDNzv4vaRqQyDEDSiKJDQK9YAR0SxjgdC6/VeBkrbllC29jczg/Ugv7l
1asdn8yQM8H3aE4Zawm13L7xrjzkDqHshwmkXyfHzAuzu0WcGxd8Y5Z7t1LAnKCn0joOATKIjIGV
EqD86yfBysqqYX9gNcYsf892HZeyXRfBIomg64Qsuxe8/qkIEcrUpe/tAVjhIrE+4u3Rny4PteEp
q9mTzneEWBmZv/kb+mzcm+yXkGaTYai+uBYfsMzRxHAai6h8Iw0D0nvPvBVefFJmkpjFLWFFzkIQ
GsI72vPiTw3IBcRnvJUB89tGcXmF8CP0aGkZ/dpKwUZf8YlPg8YSRGvOHfcHCM2IEtzG8NMwa63d
zlC/kaMIwfzf9rFVzdEXlIvwhyPk9bU6CcB9BQ9Sy4DlTtZ/JtCOaEO4LhF3gyhkQCGCz3nhSEbv
mdWJsmJl2k27v0Iq0CChNl7JZz6F5GMR5EWGJ993qXk3DhTEZS8g5JdAntj6u/saz9HFTNl08kzL
kq92HszTYZGywnbdEOjH59g0f8H/lcQRpRGzuTtDGPB9jeypuMNq3oZ5n4vVMIK+wJWGtnbFO3lB
ox523JIvXAQyUKv+ANLoJtmASvJwvHSJNLm5urpTSmfmwXJkKA7OJV+vT2WdWXNiu5R0Pb3mrSaw
Y7dEDUjMuwVlWaKAjdM6Ti1Qz8nlM4Jx9hQ+08hAZH5e3xkl1IZ/d64F9ojX9OnVmT7mhnlv7YyP
3L6rr4i8V1idzfYYE5xKYKJGe1noqN/M3Tw3hwrtsL+PcHcVDx6IHcFgUntlJZn2yBLESmpXAm0P
/QgvUhmHUMn+mknSfib6itHq13XCacNLwkOV7N5LYrssYAulsGUIJLRDyqckTgvXSsy/BVBn5a+y
ReNOraF/ptKv+sbDBr+FjOXnSah/Tr3km5MlJ5U7LoGYLSEpxX82ygdzdtvqk7axyDzNTgYApccS
hbZgh5W4+VD4/2eDjv6uHSAWmv89rwseaQYbA6dcfxPsWg6vPdiN1UmV+Oi+Oc1irOJ63zN0ddNy
PH0pPI5rig+V2lzdT9h5flq0HSr99+v24n1XBW1FZsDInr/TXSAfkJzm9ABWgKCB5/FEfMwx1car
mju3nNuV5//IMqCqwCqyWP9cXufFOhKALXHy9ZwcfVDhRsOi4vP5bD09eUQebIbHmnz7UW/4L40i
h1HJlHP7aIZiL1juqWJaZm4FHmuzmaaBN2LQ6aJQohuMaGkk0fSxxyGVZ/qx4mXZ/+l+RxwuENbS
RXvRjWLBUlzM+wRWop6B5OW58u3J3FEUZEEPRaL72pBHLvitLmZXysY7rh4M/pkOmf+b5q0nQIEW
NVnu6Jti/4dMCf5os6UfLyTYhaR5XD1i5KDrolrv7d7BBluRUMrj1gFowoXpLs+vlR82zFkJakml
T/d5OHZxczVz/orOnL2Cyr7FR38eDM/K9nnfGhbmlqsIiGymtFraZKVBeqVOSsp0JQC13xXICP0z
aLZqtGmb3SfJ5xWOGydXJ2wurvGX7RU+J6PwJW580SCLYryFlkuM2bAqvmrw2DOGz2HVBm5rumYs
ECYORo3t5U03F8ZeAzY2FuuorYW/d6J+pZ9LOjgubf4uz0wx+9Df7mbvY3KYlK67V3e3/in+V1n4
Bbe+c6LDWRqQq6y3jWsXBfHO0WBXOePIMUNTkuD3soqd/leNvpxIj/VnIMd1r2jIROFui6kdWsX4
i0vlJnkeQerc0IbKOhUajYawUUXhmqmOBNRgHmjDGadfG6nFA0Od3eXJ+PzAYvhrbbjVCuhIP42z
UY2VeC1dtzImXhvfM2IZPVLSfDc9Bq/qRoFtbSp+b+N8QP5CJ48eaNyTeJdmYdBnz07DBTToweCo
7TsIW8AhpP1gLqIlid09CldDZ2Vb3JrJpEJ8/0xBjJ8B2QUr+G34KmRKgxi8Xn7SSds5+J3+CuOX
We33HQkP2nPzxTn3Hk9ZtH22AP73pKZLbSckMfexHPjfBdHiG2OYxy9Ygoli5SUPi2sJ9I2Hehk1
6rb49Nrav+AQDQZDtPC42MCXrPrdIeVDUi3M8HOonSxWub2n8rA5HYJROheVEV+Peew9JUHsmlB0
CfsRbLWAMgccspTLNDafvLv5ljXF824GsJQC2Xz3+rNB9jltCvwfpGPeyFVZmT9Pwd1NvHZ9AtA1
GuEs3i1z03dxXkopFfNVXnRTYQlreavGXKf0+PlU6KORZ+YpIZJ2YZCLHKFrkdVDHvzyK6zewT8j
Sab8CGZCXucjHSHP+M+UMK67FoZreItwoBbqb7rzDav+zvmx4YsfF0OXAFSFHgxiS8CPtOI/JYRp
Pvyw692gFdWKU1BlWktISRGb1+c72nRRVtJsuuB0eW6JKSYhZuCIHOjYgXUHR1FlYmiBhP5bgkwo
2KgDKQbArE1yNXOOXsxsX8VFKdC/SqF9LP7lkdbc0lthLTPWfiOinluWoeKzLoKCXUH0plfcfpo5
ipbmUU4S9vkKHpzRDt7Errh7SRRN0pUyGvQTqb6GcIv+aDYmumu8aWHiJZbqPAwfMVsarA9OjrQc
jKc29F17mREl8Ub64dzuZAXX/Qw/AtstoB7NRbbslcc506/DlEMJveG7wC/6Czt4An5QwFvIPLKK
9VzECyFZFxwnsSG/ZlFkgCrlsG/B1kR3tc5tEGkE9kO55iokyLqXPDZmBAKNH1YGN/vTT5FCclIO
Zf38eyomiA57wbNqj0ybSEDF7lXeOFAc08r4nhd8093h+bCAmGL7KeTa85JCjK+fOGibEaSa+w9r
BofgsHxCtRziXuffRkCLHEo5Ze+ag/1o3S9Hb4wPZfPe8urqwe6Cm+nDRdyhJ96AWFus6Pr9Bcvw
f/mBMxTVupfLW3MZ+h9wJGFELr6mAlUfHPDk59ivPhjyeBSay36REgco2ZzeNhkQiObY7Q9KrvQr
O3vX7WenNP47j3jlDy0qztcWG3sXVazw3P7HkeSBAiSPFZHAUvuPLRVKTGDs7WMrF0XHKyg8saRi
yS8GbPcHYOWAWZEyVqmIXZWsNffGinORx1tcyZAmmd8fwSuDIy6FukM6A4ztupUcXqIs8mPIbqp+
IxwamBEPDsOjJef3FH1FSgR3UPwYHZm3FjCTamqL/A9eQXcyFj8MGEMJkH//1qPGCboFt1Uy0U31
Cm/+tWPr+9HPJnthmqIkGYNmcANCUVgbx9BYyEMA4g1J4bZb9DeRosLRbmLh21YxhAtoR3Upb2Jy
1pG0WxNjyn/nkyz50jPRiXy2xk0JAaZRZB5K2DRXtrirjkV6FH2dhPlMCgFPiRuSqEMltKJmeDpk
ci4GA6HhAYTMWsd8kFUxgkT+dsupELX5Pxx9V+Ti2MK06kWkRfuZ/JanQj5FQQh+NyZQfhs14Z8U
DgFvy2EMlxX8mT/j90OVVYszRXBD1lRfZJvbyB4qkbJPNEjN6TSoMgSkFGkvIGX/ZIVJr60qwr6f
AuX5oZzI2Uw+hJAAn+5uz+Jje6J/z62daNNjEsSke3hj1QfFDhjUy10x+erOAGTh4NZPFCPLBefA
iJBsVzW2SM8S2JKyb6wuFMOSoWu/RursQqUQ1SY+Goor1vCc/IpegqqO825z0a3dh6yKei8c7UVv
tWOOFD2EnVCtgVDJLdekDlcvlq5c4b7MGWmyWn76WmqsM+jRTmCqvjDvLdgmqi+/DngFxobdjD1M
0P5h6Ob8uZdIfXHCQ5EHPXRskxYVOkrGxFcBnjJWSEXcI4DAIi7TXulhZh1Vkeg9AkKzGZ7pDnXw
D2d/kv2BSYbDGvS0G4KheuCMFX52smARCOyeosNFBcNpwU1Qtg3t0sA/Zew9LZ9XUfADwFkEluYK
kNpSOhsf4nDRXPiH/XOFlWMPS4orsBS+5/QRjWP25uopKOuLh2tbK+7dsWiSJUg5dUH1pq0jEuOU
E89lbW8S7B1RwvhBsvZZLCQe+Iyglbee1N8Uidon+6TiDuuQZBkKCbWop+Zccl58iMlQLR2BJNhv
fxpBd8jaToTDsx09i1IQ8Xwp/yNQhv4eOizdRvDAxJbAq9tRM6UOZspp3hdaiR2zsTAJy9NvGXSK
7NPSRQglHKHEOcFQ/iggDJyFAJ8qbq7VeUuHxd8GF7UjmtYL1H6Ggy2ABeejRkx+Z0WVujmPR2nJ
gzo0eTQmzc//IbuSx+j4KSHnYdWKYb47Wy8HvzQ+MWd3TwH/1blX35YvK3Fo5zqQxsdSVJrhcelq
bIyP9NPRYf3RtP+Mj++2je9XTGBZZzYxuG/QqAQA8QSuA0NiOLOHZGc4r1kc5WPOL8/PPqDRkN/U
VHmzfRpjSaECV+rc6jFZwgWWFH3PeYGrPWvFLVIvBaUGsdqw45T2laJT5ajkhzPY0Hi7s9S0xpvS
VjYpTs02tYQiVU0jTU2SIQzXV/d4h62ezeKb3iWuSG6jJnergW70HVgIbJw04NOT6kKfBZuKXIuS
sfHHyyRVcqpj+Jii9ZgF0qU4QtgZZ6GfUBynFRg5z7op+CLcpy8AgY/InQUqowLEDF0ayxjQ2Qre
6wMZiXYmrNCKuoLbLAuJzil+xjsZhzRrtcYUxwA3UMzftUGGsCaKLonDhAXXUIyScy13uefsik2b
xARPQ3m7xuQxE6rXO3B3mXcB1mm6dgCQE371EOlzHohNo6nAvl4w02XDK6tm9k8EA7b4NIRPGSwA
n3u7D1UDZdAB6VHTX/KfTM9DS2XeC5hUZZNrfmwUdKnBg0Fo+u+zDZQH5/UWafMK01Co3nVZzNip
zycqZodCC+wbQ4T90iQbooyhhaoFM+XSqLBiNUeZp7qif+XTvS+LPbrTx+QfsVZp89MKH6vX9j5I
2aRkhWs0ri4zu+Gl+AtILZMONgUHaX/FFJQ0mkLsMy2J9a8CEuu4BEIfC1C7gn76kj58quVAM7em
Rhl+QBQdm0VnofFhPMfY/XJq5ZKLtFsmKxVne2BYp1sX0OJAy/zkLVtx4brWhokzRdsKeoL9BXDm
/PsMuR78jPldlSWCc0eWCvtgiH9nDNLSc2B/7NZm2+h2b6PpFwopszFCo/PXtwSF3PmaGobhI2pP
R5rVK7bq+b4UEnYmU7jU+QlSMVzn8rtqyQg8AaD2AhJxM9890YOHZDd1ErdeGqGGId/58plz324q
Y0w/BV1A83KjKkGF0/EOzah6pttQ+syvCoGfDqZHlaz9i8TDvONb9c1Mzi/BLO8PfCzk0zvmdIZn
08bSi6Oyi+GgKJkP8dhky8mnNcRSegy/Ds8s74ElLawxm4ety6KrHbGts+F1WaDWOcDghEKa1S8l
RoaXaxSyJZCHgQmqFov+sKd8pWtnnpl6tQiAtLBrY4Lg1+L68qyGz77rV8Ybcxb6AiA4V1Ack1/m
UGHoOErL2LTU9WsbyT8SyMSDNBIvKEOVtCSU476iRFGnfKtqwoK6Z5b26HQophzP5TNQqIK2eoIs
UhT4t48QS3Qb2Z7nma6pHL+PQSIy/K+XiiSYMOOA1ODyVNagZys5KYN/GV+I8WAVr0YaK5QgU563
VUtHb54fDaGz8S12BfbUC9b/90NmIBf9jYUBoGP2P/FiYr9ts787W7bYbL7/9IqkN0BkUvmsE2Ii
U6Sh/rsMCKSFtxft3YEAebLWT+UJvdOs8WGAJEzv0jSV35pdyGlVypus3z+5rtPSH140gJuzbQqe
7FtzzO0vB/9WdkSGOk/b/5g98eU/7bz/6MjX//gB/JZRX+9mpkW7OzNMdgUvs4X2WCILuaaJhYfp
2wtaKSzNlacxHHfUl35olY8jqU1xVTE+PB0JWkKXwSi/VyNLiprP3bJ7FrIScT6aeWLG1iBwTY4/
SJEYarEtem22m5QVmp1BXxIhVqJ0+76b1qw+2tBcOy4+NHH2SXtwKi1vLl2WZUNdkOp0/Qff260c
duop1+0Qd6+ek7zZq+PESZbUxh+wf0NPQbfxTGxkrOWBXugD7ZoeA2ENFpxCPgNiL2s4Sov3+9Qj
NI4RuW9dqTj9w6BOX9FDJYQalq/LGpxTyM+PtooRDkeLkd/9w8+H299viMfkcqtGqrAwrfVk0t5E
wx4BlhpgX+jTnCFnY1XfTN6rdvn3mk0uzjbN4l8XuNGPQTTzqJmkQGUIeousUUKKAR2FVlXeX2jP
ESfBlvb8Jg9iHzaGjk+vNb682m36u6pbp4syZZLlDKr2PDt26ayeXsx+WrBbruLj+wx7Fem1VVuu
KxUC1qa47a805p3i5ZEFW0lICUm7lBe0iHqifDib7GmL3OxBjvFUYeDfo+e3lKyno5v1ETvWmV9U
YH7+PogepC4Ihe+ijuQl73J+oox/YrqsdAqfHHmRO8VREoDvUEWgUeWMTOmXSUwgVJsjJwfGmYCw
q0IXTQBHiz3aQEqGlhg83IV0fFhttNcSTtwXw7/FnTabbrUgabBBugD5J2xp/d3WLyvB8Rjn5fGq
ZaCByCzHADaERUq+xtiFXe3nAo7f/N6ufKkV7tX/AbizO2KAHY2+7wZiuhWWVL+uaLuPO61DmaYn
sFWYSGYntG5IrPv/pjDZHZB9OtG3rNzcroqixI23aOT1Fa3KYyFDPIaPF96cquf8JA5xqQ/WxiY5
opfnSYHLAjDyK4ZvR/33W3VJnYYU1X3J6eg7kHCTpaf7JmL6rfJSaW1XHUUFPfl5Dne+RHXxHSUI
Vny4jvHw5e4dlFnzLeuPAujNPsfwMb/UKsu6FQVDvmwnm1zEnj/9HEczA1yEd7LWffdGmJTjx0cm
UG6CZzsFXg6PsIOh/Dg12HeH2NmYcghAqvrUxk83Ruk/r1Y7+OFH6snOzfElf1OJyYqkDVq9qNkn
9dw1rmrN4j7FcKJRCZPkOMDOdBxkt+AYB68xEXOTulLg0ffZM1x/LGN3iGJF9XczdDq+WHurBw83
y6LgO//8PI/Zadywo05hutCOdL8oUU0U95h7m1kiRcwENe/0LefWM1+EyPQ1boTWE/W43QA7A1ZI
wlMbKBrSSRYH219blKFbSGquQ23X0Zc53s/DvaSGPSiSD2THZu3OP1UR8h6KOyXaSX1iQGM9+LFM
aqTlBloUMbhgUi+3plyRV5VoYV9BPaREfjxUG4oS2HxJUMZKyYSZuEzmeVGdzkXxVz90GSZ26wu9
GnrZ6s6QlaPK0ZMgps11YxcbDlMMNTTVMfRETO3eumojVzwGdq3AK7fCA+RpPGrUJ2Tb+pDneP00
ApLrEalcu3jBGzw9XmPmnSV/o9vxRjsbvPqAPFS1vl/fzgtcF+r0bHO7y8io544fDLlwGUhjbUgm
Yn/9oHWS7DFTGb+kheSQDLaFndKVbNMp4BMD0+ouVwy0llDR0UAW7tTVpzz3Ig2MeAKpbLK0Hn09
I8t0sV+7ntme7WrPww1GIZjz++U+TewgbllxA/guS5h3RKlB7zF3Vql6iFx8NCWTnFjbVj6nUoAn
bAFhEhP5MiEm2oSwYkHUFsMKe51RIVlX2Z753MEV8L99kLFAIxtvNxn/VAs2Xirzq601M6AvRAT/
TIgXLVNVQ5Al5+F9t1+74NhdAFGuF2NwvVfAOp9QzECYMuN+nQh8WU2tlU7wwQNvsxEwf5kdAHY6
7WfuPoePeA1d8iBQRtOG4DDwY6J2lQVLZAqkj2s0Vo1cFZefwV8vJPAPUTC7Z5oq5PKiMrG9u4xl
3bIJ3eBgimEDNCW4A7/4fRDoDVnYt0PnTcsdyQTOvHCI1YC6aUKu0IrWtW35q76S1u7s9ovXwRcI
nSIA+klZ6QyBiSpzz9KMSCrkYNz+axC1ovvndc8uIkusv4BlH5opjmWEfju5CDpM4PGiTuG0jm8c
QSTKYSnG/vI85viCSpT0D246dGl/d7H7JXBlmrUu75u3043fJstgk75J5yRqB5BGw1cWh2WOmhI8
YtEGAlbs//sx7rZ7FQVTDYpIlqpajIm907kKz+8qlUyVkT7RXcGaqmQyV0Fy+2UkCnI4eIiOor3o
R/GmUGi1tU6pGQuWhwQbhLEECl3mAnwaMdkm6GCUkP56DxVXllwRIhp/nC2B561ActfGGdvi0XOL
3PIJS6ui2akoOajkLtrnyubKty4lmIc35w37lB6hh7idzTqkTIiNcuqHT0GUjBShLuC313eHszcW
HN/Wrnws73rvtI7KkLxTt+TMbvm7p+SX+hLqA7on4mTiwP3mNDCUxYqx7JUfhWgfCbK0wI8C2YIR
KT12udnoxGVu3kNNa6+9CvixAtqhvoRXalPhe0ViV4cgnn7drM2mFGXr1l0+WF6IOwgC4JK/04Ka
qnyQe16L/b9LnSlN7359NO+XXsW41TsALVt34oJzKcrx3ZX4aJceEPx8zizXD48yhDrt+/RQs+UH
+M8PTUQgpxH29D/RMLFM5IocwF3h/yC9h3C3XZiE7CvWv4AChvmxqCXZKT7BbZNMfV1pojDBNpxg
XUk5tc2ijHl8GDjcCyqKfh66wC+tUrzpv4sLx36Yp3ly4wABkQJfvjTk3zh2ngsxcmNafUKg1+hE
6XGMtKA6AWPTNinkpiGTPrSk4da7ss9Oh3G4JumG35po1c9yGYQsljML24n8qkM7eLI7wfF+TW2f
UwUWNJDNuMYQpk3GtSgMzMKL8mSXhxFhy28ZLtOlVOd8Isbw3zbsk+yBbiQwtiE6zR3RnAqhwAFI
/r9xWI08ymueXX1SMocAd3LiW0Be9eSM6UWaAQr/CzvCXM+WLILIjKeOE1c9cVV1X806kbRJqtFt
1G4i0oBy+iz/n+gDDUtWL22wdBRcaFIgJGplcsfOQCBYuaf2ufMW8HMXLU0mGq6qTLawI55bWdD5
9gdcT00mclo+RwkJcmZndO1pgx7PCnUBuangF0brp1IWfwLRK6Bqmzu+xVl0BTHtzRpPNC3GamUt
jo8rPPxvX4VAkzZavk0Tj1Rvua/7RRbMq4wNZ+AyZVWZ01Lo6uz2aK05Za87EpZa1sRXZwhuBq7X
C7LjB1mpf0zmhR/MWkHRPnHI5i5Lxx+Jj01gSiqYIP+TjVmpDMNJxV88Xu8yY7qsFpKMopI7IQkv
LhpCCbNVCc6cR/2pS1b65KW/DZ7oOQaV+NMAVbqRpB21n3bfqoFRnkqRrFwTPQL7HXqbbfaorcBE
VOou4j+Y4WRZm+oEN7WycSAka0IPw3j4+2yXXqOIZHTP26MUclGsb33sd1vpJqJAEKgTrQ+mPqh/
muiX3KVjqumU9YhIKBAqvU/d16eUYujyWfiYi2B6mWx4QdjxDqMd884GihIEQ/ri9GnkkafMEe2i
jGFsWhtJIm8aYRVxKpd7OvYicusjblyzwppCzDVDafxE4iCpztvib03Nad1XDvMixGrS72VsSqMO
uK4/pd/eWoii2oRyKA2c5pt/5RICaI0HXgJG6Csd55YqdTdeGxgmoocXXrKeTdMLTvxQOjaaS467
7lhgQYhnqMaoOEEjCRt7iCWdU8W34mdWi+6xgcN1t7ORplKm6graVGpeHtu9X+P8DULx4h0+Famu
L7cnyiYHsFqaGXpjJVY3XafAW/GrqlRXadeyqWUq2Lf+RpgiBoOo+l/zUxC3T/ac2QjpclmwAfrL
bD9r2/6z74uI/3660KKvN03tG9eSRi3wPMpE1upndLXOCuEp4zaHgLuB7Gv8assLXmBgofuVH/eL
rSL5vbyrzTNrm0NJMoHfboMGGFnbuFkb07sebwHpNfzMKqSodFA0iUnqVyajlNA4bZ/WTAIS9XLX
wH7/kktWJHwIXI8/MUpk3exUebeeSF7vR1PIX81sl53CGjA90cWX8LImVuzqm1BBviCbDH4n3r5J
53reOg15OODXnwkhQbeVJKJByGMoCjmcbGr43kaUChDBjo51Vr+rcGp7GsqgJYP4irzrSO2lYYWs
yM1zysgkKlJbzlksSPT84mRcMXfT8/HAndkV9Y/rOqvgYVShJDj9vXSyAU4ooqf9sDBiZ7Azujpd
Z4MsKhk7UrXOHWWqdE2Nd3RDxnknMVyMjJ9qQEYIXUoy6/oxELi4/tWphZ3WPotBdLD4DqmvRAfg
YOW4nPu93Cw5oFHr7r4qkBj9BVOrPLgAHLjwaWayLfT/ZY6MUhx7iJ2XrsIC7OqyqBUX6Ie/4Nwh
q9qX7TxE9NcDgSOVcv5yCPiT1E+lxXMfLPiMdW5ybC7YJPBA76vH4I6nzbmnViG+8cOMTFWO/HBP
hJj9PmWrwczB5MbKJg8TXIOyfuHGgSjpz/8tPCgz2DPlgyZGgVpNgoDH4neVX6E67ZckIUHqJQru
GcBoC6QseQ6Y3t3wJWECcnjeGWXlIY+mbGMKzdOm2HeDgcSYtzAEUZaffxn3Dp2CS0wJyPCWY2r0
5Lq24qSA+5vqYDSvNz8cIlKMI4rgrkIujPCwXcuCMTfu2J6gDbFnmjU5bKbXB192mNwpXCtGHrUQ
dgbEIg+dHy95gshcZdJjFLc1HpNa+02T1n26EkIIZxe+oHBoFTvQwPG/fGMxSL9PQNfrYfuxtK6b
pFagtVTMZI1ZYdfEqucONCE/mdXNMDisrXUxvghIvU2uFXpKME50vsL0VB9erPZbFz/yZZc2/KFM
nStfC/TN21auc4ouaczncvnzwNdKCWnpLb7pPrJ0iaZQIbdP9CGM7W7YdttwOJSuZP6sKJLHoQZv
z0ouO6Xcbpr93lE6E87aJSJyQm/I+wFmBQEyADwqKN/U1iIcvpDwaTCmo6E2QJgWfLYZlLPdm1Kq
K123O+a60rOQ02szaKpGOhVQ6vpgiE7DnHY/ioj+XVs3voQ60cEW10bXbmssHiQODIo7v864J/kG
8seJ8kcidvUB5Dzo3tXYrui42Cs2w4CMBorBA40h2yl53ZIlclX5g/VJrIBc9FqXZShac3DTs4bu
61HLDoaErJqbcRvBnCx08ROSPKVgCjs4mR4VTf6p13afhsMzo83J3aoIknCTjPdvuWQnlQcOUSUG
bBAewYsP/aum5lQTBLRMy5KSbfaTyDSojEiRaukEoopB91GKUeU7UBBZug9yldeX0rHsJpoKQI7x
aAbXINp4atoGkvAYUq9nk13BaoBrpANmns0gDH74gSmMewywodtC+nKfhQXeNMLKl0DpKdGMIBIi
bePmNU35OgQo/igl9AWfQN919lK5bN5wDoP8gIHZCW2X+Wwv2rqlYfLSjOPaLB3wHzLSZ02Ye9pP
J2Hjz7K2inHTMApeY8/Vt+t/zVvFf7QKRCHslNm6ndsfeLvWFN7Kenw9DVuYXaIrisXbdZFXCNfy
61eWYV7yYiuGqJsWwvSC07TUtZzaDt61R/SIdIsin0u047tX8BH+QRYbp370H1lgPgTklCvySR+6
wN6kSP0ppKOn5am6LE1wTxB2qqybxtOtHyVePYvkWBvD7s1tEpRpIOS+W/mEBsygz12FTJnDAk5Q
kECtaK7ACAQzHUGKTCRpTrd6z427c3utB712CbEcbEh0oTfVJdY+Aq1ILq+6EOGzAinlN04lYk+M
v+FU8KRRuIBa32X0bFwetueiOP2F6WzqEdpxuhiaoJrJ1OhjyQ7QijhPqrd7KsouGUU8vWOAHvYu
rTPawaENk8u/JgEV7WIG48Vkz051CuP5w1wTLc2nHFi/BpXTh+yaqEJL0RZiUREb1jvnGLgR7bLH
Pst+LP7XNzCck1OKPlYWdeXGAvDgD0SdW27ikkGN5HtLQIuPZ8Yj7/nMrT+OaUsS+gSCGEtuiooW
F5K2+FY9oSwzxmiqEvurKHGKufKFQEnBGaya4cXWFHZftiVqtuJdabiJzDcJViUutVO4tBkiK0/3
s5Olu2R3Ar7gXFx1a9r2J+3dV5/6OXRQBW58P7wSerD1o8HtcKXBOxZo/s06eRXqTeySVfrFqjaB
cc2CcKEgHTUzucnEIm/xz+HtNET1j7HJv0VkStMmY6yxhvL0Nl/jF+hEqaFv4X9k4C1F+aPP/Vny
BqBjx3Ny5er28oNhT5r5MW+fShn3TPS56uTQhxnh7iKeCecFfcOpeGg0JBaF74l6Kmr4enmengur
s3rpjzaLXTUxENzjuE0CwjCLSrs8C42mluVfAeknKVYUtfOyqgfK8FOs5aIADdKPX6iAhUh3jOdS
PR6g5HBF1QehBbss8j5ojo8JSQev2ON8pUiATaFqeIOdH2LGXkrY4MmzrVzVe2/kkIH4lbO3q5i6
IgwvBGcHd1qOPMegQ563xgL7xW02oxf2bFRrWZ0xlRtw8znHAC512jH6wI+YXCElCnwUGQW4FPcq
EabTOL3Ah1YaMxSFhVn5G9gz8NGq9Z4jGEuiw3nJVEWlUUwNrmCMJccuKagGIBBDCwt7ZQacWQxT
C3h9QX31HY1fTuqdnfRcTWss757Hds70scJvBqVzq76C0Vld6LapymoERZaOsvwWVNyUAbxSClb3
7MAZEwqA6awzR1/L7Qeaxz8IV65QRWYVqFME3zyVH18iSeCL2mHB+N2YTTVbsYwuhVQ8Ih2ntHYw
8V45LgMs+0IjJZC26jJjJzUV+NCCojMZdOyJm8JHurR4ABAORbkd/0SwL55SVCnYDmssMA7RZ0Va
CyoUPdU1WrOvrEjp++CDMfdH0+cpvLY5Hs9HcrVv2McKa2nZhgk7cHERCawL1EN36cuQV9FOO8JD
qCliwiZapP7P9Jt8N5BOYoQVBC6eksvFH4J1etbcGVIf+Iopg+hM+Hb4IEun/io6Hg3fK7FL+6h4
zqVFjOeFHz8g3zN+Vxmh8ZzFJVQ5uERsYIQSUNB7/kfF5rS8BlS51glfG/ZXlpaSz+2Y9s/OBq/f
tfY/uYWuIPzKhTjDmfOVU6ck34iKuYhg5iBXEXiNg7N08ioTZAtze3y/VLjgsufyFmYlhCKOuxgY
zsqzw4FLrW7hPgGRJ7hx09BXiUqYdIM7pMQMapnfrYveXf7bOQ72FnIZowKUdMpwDXXgyv7GSzkM
sNqdYaWhClmNfRxisI9YB8mRs8NBadV8ou52z0uTROm49PNEvmy0wX/n5BKuCBG/QUzxxgDgyaJW
iGEAbvh3Bugdnq5VhZJU/UYeO9/YFPU/M3EIrG7yk0eQ6s934izfJofmu03HxaMG9T7IfAQsyRhk
c8FNbyz0klaIEbcnxU/cEeK1HXfhS/EA6R2jB0nCDs+cuWU6nbDYHCaQjqhmlqXN4lJAk+eYoYBf
Pf5ESNfdrCWRqzBu5VFlANZjKt09fL4O3L1D8Oce9gBxOfbQc6MTCiBW28XgIUUAbwGynXOiPC0u
/CeC+z2WJH3KGfp/0hFw30elOkhr50dM6Kqqm0F5/2L6O/1QuPxrrmYbiJ+5geXsThySjEb8Aa2L
WD7OxuQrwAkXqRJLbWEwlQ7b17+TPFpnfOwN8g2h5K+p20iFP8polp9pddnBlEFXHg156eliU+qR
V4fUJGHnVlb0RpimfHFOj0tvqv6WxI7gWGyUupxk7N4uMQMIKy8/SEsZBgf0EudAAdpvtUfX0TWB
rgGMErHato2nngMN/pSp1mMvMdrgbVLx6ivEA5NfEw6CMTUbQahS+6RIs8HFEAOUsFuLrr9f3EeD
074Hboq3OQCHPT5ggy9W60ADJIK9LslLeIPL4xm3pOjQv4TjkSCwwVuTOSyXwN1JaY7K3aAq3Q8D
GTN5sPpJGgW00VOPP6KUFmxCjQxBmvO8jk88r3jJaOWDcUZu8n57a92m4FZFAJjQjWa7933uINCB
B/4UuMX6lAAU8kvvLFWi19MRMVgTAeF8ooUgm8JBFmZzXAC+hPtr9EKvEZ+Exewhekh7c2HYhAhf
kWBRCG5GpqvUepobd193wbnUCmSHcBhsoqhyLqjv931tbCmdWPdhJ4AHRaSy2EOJxq2d/8uBAG+H
v4Hv2Uy8SxcCPqlCq/0tiV5/fXyuPYXPg0kGy/0ePevB+g6k1i0XOMUap63yIWhWX28n0yQa+u4X
C1pW0H5pbpWfFSyJY5GQwmv37Zj6SKBoavB4GFFIkTq4vwTwk2uxRqDHNrdW2qEBX3L+qU2OGG4g
9+11VeZ1KrglZj4FoVZv/ZSpY8xZyiH2MwqfmM5eiet8+ty9WuycTj+I2MTX8j6si8d1Tp2RQ830
wutUWKDSwfA/nq96LEn4adFwkDHhKrhHg6j7hm4Ev8pruw84z/2PIJBcF0oc00PJDECS/UZKcwd6
tF1ciVS1dGNPnpPlIaJ5aAhXBKwRRenF9jRPta8+L473KXrDlJa6JpS2C/JApJsyDrWnEwBsbt1Q
qAYo41IvTw8O9C3mPbyuy7nb5p/CX4E++mtNbRtLJuIN4dRxigODoIQQ47JWSTpZzUlZtIm9nwUd
0nowv9Cm70niwNHMBuE5pRBsMuvFEzFuefRU0vXQiYnKTHibG7oPNlAcDIGj16OfbqiT1T1cxvZw
+hQUJ/x3DHvEn2fie4mC7BbXstoZQ0V9CTKVOEK8KQ4WqLbnZx47Lzz0SfFjEYu3Aez1ZMQVBvIX
LEj9L04erX3vlW65PQy9My0V5HOe9Grp+mPYTacnRM0GKwV5cVe3jir8XyLm1hUqNXtgskbxsdYR
3KuVvJviCufsHFMnv8qj+yBqscpXhixDbxiV0nEze0L/zxZJdJQuw7BUdA5drZjAf1S5YClah6HP
W2sfs5dR1OuriK+Q5Ko2obK9LTXrRdX8brTICCMgAFEpAfTgmfPDqu1smQ42vlwqonGdl/ymhQtG
NZx2bZcdAsaiWSHbAoOssGmxrzupS3n0FL7l4vC8e9vugdPBiNWl5+cqpMt67VdAaiwYOqbk6YlX
RETUFreTxNy5nhFuaXCGXCJ/Oc88hOo/G0C83ThSiuC0ebj9D4U1EX9hU/A0q1160dz5+YKuZfw/
FnyeyVzotTvgyugVkpnna4M1Ju4G8L5ezZQzI/TD9K5zGDf+NejuGk/40dEcSjILyGv99HTABYIf
qKbdAqhJ9z7JVitENPsjelt9oSHvFruoJOqDh37SoEk8g544kp7Kk+/TGUI6QZlqlyPHNYsa5E5w
1Iqul3eDIEZraouDUROoKhHIC9nkaXt4OOE08hQIaFK8TDrUK7AsYK8gPsedw9bXkaDWgbkxDzRz
ncYKIkhFLMK5YpxCLhXwuzhqldmjPE4wo/kAJYJUSAElyDeqe5z0nmvFZ8Te97K186HgGf3o2m5B
exMyldl0TLX8MMOjnNcf4FKIN/5ITBzsbVzwhXdZsjYWBCQoOuJMjX5+zut3CyQ3DEW+3e4aBCO2
gVdO51fouAyivDX/IYuaLY38wjZktcoRmAbTJJDKtG5c5x+aQcjU9m/mLGhD7uzExt8fvtY0+5Vs
b/Ffu+sgVNbnMc/DobpUzzhbN4fNyM6kUJSLw3Kxgq1Mn/+9s57s0v+XKeGg2dl0iybOOh/zY8Dk
5f609sXlFx/DM4/uhl73SDOWhBI4Sia1GSfjJWA4Vm4ucsIxFTVf0UUToKM6IDxxxuEm04e6UqQw
s6Gxclh+5xojSQ4F6/tlFkuMQc9uNpvs8SgGz4IJvjticOC8P0kSNoHd9zoAE/sIqugmdrk3YY4u
VC0D93UMwf4h2/U0eujTJzCGVfopZ0M8deBwPuN+CYaYO5DxNsSS+qH3+hJ0vUPPiVrnE358BZEr
U5tUju/71qwFGBPlE67m29lDoEomCn3rvRx3+jP3HTJojtCrxE86xy6DAQb0LfKmag2HgucGj0wg
4/F8ZyBHhGHE9EegQweeAWupdbFDshkefC6T22HubktKuVWSVXyr85EvB74flkPESZyfvciW8U3E
uiz3+WCQUQFskhevaPm+0EX5SG9HMoaj0rPt8IGbClPie9sO9j34IVy4xYGqR5fFviZgwWnzEsqq
0nHGzq4VCVg1WNWCFerpiIs1SBB+sa56oE6cIN5DRAfmO9iflhVBcz4tTnpska/E+WtMUxoeOquC
mcHCMO8rtM+0uHTft3DfeWcyOYpmViIYdRQzU1sxPmiY0/46xM7i9vIfuD5aPqwoINHXi36di7vj
+zfAljKDtm/QZqykWusfE4kG42eWCSoIrDOjHmHHWeOCSunUrUhiJJbX71us8YgIXu6TTKsYPPQx
T8QhR76HSlN0tcXVz7AtMdlZdh9G2SElOvGPxOFzMIxo9+4NAbOyYI7r2TD2fzNTklTVNIUDJUj7
F8pi3wLFL4/BXpjPColq0n3bFcN2AwW44uh5b0/oSs9gin2RvHLDTqgKxZ0z3KfyRt2WQpIlttju
nuFKv6oHGTwStqcafPKS/6rYWPsl4mHY2fkEoQS5nUovx+gfE77KZLTh988wHKxRv0u6uQQkQWuO
LvTZ7V50XIOVOEImT6uu/qHgyp9nKy8yCEiF1/AI5+pVmCwWecbbV5CdSWUeGhq3wlH2MgleZDSt
x5hVAK6PBxOntZxon1HkuwPPLDGiABl6SdRJYM96pxZQStmcFHTiG+IXkLjr9PipoHwhL8k94HoW
EZ1bjwG6S4bhpC0XGLKUfHfizKCl4wcIdOWKlmq4F9LfHmgW/yYJsatW9nMNejvrjiuMgPAK5J9G
1fnkLS9fHKH3anwzse3rspV30En+SR5MAnFlxP4cxZD2991puCqJ8yNklLvzjTa6z89oVOAy6D46
E8ETDwDqqjycFxpO85sG2h/My2Rcgsu1JMgHoqK0g2FVNffHCEwGFrWiNfYoS0avNNTR92oxHChJ
m/ufApNZ7vAB6anrdae6CQDJ4bNTqRUd1qmIYX199SQGMg5JnOqBGu+HUYtt55LjQSjtsxuDVT8n
8N1X+Tr1RjQOEWdC7LkOUvmLvRPPzknfMQnO++CzggtGAy0Fq8ASyNpfjTPzYxHV9QoZRqrjlbRP
TjrmmdzLB4WPeLOYgF7SU+FZs32RinyB3QJoTzceX74g1SEOhaMlF25h4+BB5P0vBonkPX65O9kE
0ybigoNE+80mW14kIfyBhDYqLCWFWOjxCa9zTJMzc7by+pJ989FhYI9F3fjqquLOamm+lFpUxdZw
aUGOlDw7U4nEXc8jGaQifksoJsbwjlp3ssnYqyLMHiZmxeWRGi0AsYoIxK7LQTdJdnwEuXiq2mwA
TKtvWZ/EKF0DM5e2ws8ZkBneRZPf3Z/WsesbXmVtBj2uj4xwaPSgjDpX5ZU13A2h+Fzf5/qz0c+v
OIz1qpYcIy6fJAHFqlGdHQq6KTp3K/zG8t+lk7iSWXUyAyTcnR2J8sGQIlb/p+T6KlfpJpX0xnfT
iF+pBJhz3dIXImF7JX4m2BivizRgvOXKJ8ZtITSWagANLv2/xwSEwSfRMjxcLdI1OjgdL3xmQlt3
jp/9dIDb9qxFJ9WJVtQi6u4WW6H8wmwQ+PIFtSH5j0Z7GKWRoZHlwwtrhqeDZRV5ouzYs6tyGJ5r
BG6ih6wQdQ7Z+0w5zhQrLN36DN68/jP1cWfFfd/IDUf5aOpIsxJ1edNDrn9B8QmRFZRwT4tO547n
DQx9HyBOUK+Rcc6EITpeT8q1PlrpLl2AMQTuk6CtlfFFV3gkRJxxF92xaMNNvGd189PsQH55W7/e
mxz5Mw17VKmzYoEjGxl4Xf3NgaAmJXvZCyACiQasbTxxZLZ9uN1s8LFv7JOFLPcsGE6qGStleb5S
5w/9pBtb1XRtPGF+jLToDN7RGuKPUsJSFsPGr2Qm4aKZZgd2dtbz2j7xqM+6+x89dpKTLD93e4d+
XrBi6DgDHEuhNZPsFPWtoNYbUSYjHxUmfQtzoSVTNW1HJsGnAqX6bDn+Wy5g39uNyDOamHl56DHb
GJknBfP68NYZSuAi9mOFn0yg4ZDxInw+ReqI4kKu7i52imrWViOf6Oh2nzo964SA3J9DWrPc6yui
zG5QIzo08iLz4x9UnIOq4W9Zm/m4DBYKd5lbJeRcYeSyq401Wza9mBuUitQvyv84kxMpg4cCnqbu
iJ2RdmMnl1kSqngQh61LYyI/CPsfzJiCkDXexCUsNWoGCwJ3ZMOsA3GSiyiWZY5/hL/KGsH6Ha6E
DBZJl7zqEbDlj1kzVmbk9mh4d7L7NiXGT5HK9jBokaYat/JRq6P6aj84LcuKKQm9sPtIkbYLFwgF
FyPXKyFDBB6yOxUgc13YP6ZZbAFgY7P87BtdB7zaocxd+0WDhIq/BhmMFpG+cMu/KQqUz0jAQZcg
YSXvzLrynm9shUU7W0ltFnoHp4XccEwUHw03Ha8MisB/+kkXBd12dNoepwxVzeeIW4LMqgy8oPO3
sAPNX4UT93137m5v5SA0xWtNwk4IWgq3e2Nosw4WBmfaCLRlrCQW8RD7i+nDs4C11+G9ysSmcovi
sF8wWrZKLJ+hmUxRwxbBXVqtfXq/0l5L282eTsoVWHBlaQZPziB7sMzphLVKMauwQFLEOXZbGGi7
aqVk5KOKM80O0X6lRrBIjYHrpAVO7VOsytfhJn/AWCjbBNHecxLahtavhYKWYaBQTvPH32gECWid
c8pXddCo901/Ebfx4Hl3QdKaIL7N/GrNTe8JBdfzLU+5TZwdfr1yFPGB3vdzulIR3tzWu9NLnxvQ
/C4/IdY6qRGL+SMv4CWicV3LgOmnOhz2i+eAzJuSOpRXCKC4vTafwFGCrKedSLAt3qqyMiVtW0/X
Q16UgoEGFs+9i93/ChnBr/32onW3y8gLnnqUmwBIf1/KdYkkRdpo6xRRW8ysYiQKWczUMpCqe9hX
APdgH45q0faJ5oIejA1YGR1g2iB/fkTtkrqyDAJ4GV6vwcTrXlk6COAbX+DKYwW+iVrZyHAWMghc
wBAMzfrI1wzxAd5fimf5x+Bf1eawfaOvOC4LWXn5EgFbfrReRLr6m0UV9RHMnBH5wP6C9ZjGaMRL
B1lp3Hf0cimhON9CxHjnU+1hvDCshicrPdPO4Xh9UFSFKjldKD6gBNCiTK6BO5Bx3NMpyirL05VC
BLY05AjE3XviKxzcXQOcAe2i/56X9w/Nf7doTsT5NYcs3/9kteJZ5lfHVwxIiUb/naTOrvrv//ih
JBr/J32Tyh84+9cSxT5jskpMMPRgcLNntgy+AGGdVT6+BdCxvHDZOr5KqqSihNBmYrinIdbpIn8Q
DpNGd3OTj6IsjJI5VBuNUaIOG7rw7UUln+NJdfOpdnksunA9WoBzAvnjQCBkx1/yXQNj2KdtJTsK
GgFjyochg6PxdJFqZbgsXkquaKD+Id7+jmcDfizO0tScDlXpnEDQiBzAsatlHo554ffqWuu84VIi
6hAn6otDG4YL93eRNYJ6hYKVBe6tQCF3lTbBLtaChvH3ZLaJhfRoud1aXLTOsFV14gaA3mHLTVZs
dkX3p3uOTimHnw5IzSE29VkkehPr1zJf1z1qP7ex24i5znrRGW/GOhvZvkHVMdoar+TE3r/RGee4
RJ0dML3FdHCrMxgn7R5B8rz/GIsgRQLLdRfIntv8pSj8dbFbwFPjfODrJmmMS4HM2tzcbRQhfO3V
5leG/6Y5GjfpJ/JmAAnwvZv5c2CdaGpzJwutlA3Yho5mKUMtic6c8rHu9++RucnAmmoKVtMzYcyw
LgoGNHCbi0AFfBfW/iViiA7kK5xt87Gd5uyyYqI2ib6c4wwwC8EarXs7a/57YXGHiKVWqM6UJIym
7kg+hUJ0XMfcWvkd0SwM6mR8xGz5hhe84sPq9/ejEdHk2vyc9blK7UyP+XOdl5W7NMMru6WtDF8r
pLN+Y7mCgTli21FoxmmkvFBFpudWN+o5H0iMOltoEoLb2GPXDPfPHYLt++S5M2UnomRr8H7I5FzT
5KSvLqgcZl2fT1bab3jPLIq92E6SV7ZLmeDReCvgzJC+hOSjUYKzDrAlxYTMlxs+cHAgR9w4pupu
HKoDDTQ4VHq0Hcvo8oyqZGGIQzmlBVxnPszRHYonRDK2+E6j9dPS/EkTynMgae/reiwJNMQaLT2q
sYsPPkBfv45+MBVkmylsGw/FGcXZOgvzproU+Lphv5lXIiN/kCddiK8SKToNkiYQyF71yb1Gg67E
PXIYxb1AsUeqm+fSUH24A4RKaDDY/h86e8x5Mz1iwZZTtNgXDVPP7/2CiliwyU1omoWSrNDBbMUF
C2BD2e4BkuUrLnTG3I9DSslkJs1MpSEZlsnjIDXFLfAzXCPrBSmGjm5t27NMWvPCJH59X9DSjvjU
WoQzA7gvLjsKZ1s9DSQen11H7Yf7yjbcdY+arZn2xwHC3xKoDjA0H5OIOW6u/d0+GuLFuLmRxXZM
pQLm5vzlzJgn9CPXPYIWbTBUnXCfuNWaHSoY0DgxxIepH56pQQLSQp46B7zLiOceBCI4fLYCvaKZ
5s4xKj6qyxcqMKYUdwr0h4lywMZpYa5kIO7AP1d/Zmv+qoGbaz8oExDuIF/Vpk2TSA70n4wquutY
f/vCQrJoK3NsbpSkjTwo0DRBjcj3nkRYkEienvj/WrLjhrKMdvkpLmwlZF2lgxMddkesKBlauwRr
4suzRqhjmg/mNgYkFpoFXxH00s5qL0nR/KS/HyWSa8ZN8W+qO5PGWVbYKqbqKWpMPQ8JcLHN3irh
4tfvsYUTYorSSf1P4dxO0JZe3tP+qgDt2Et1ACLWVqoiuMgWbiAF+Zrt5hUxQ8nMvQ7So93Mz4CA
SqcDS8VOcUp4lHn436slVYMJHQNmgJh/QqC0NGzhHPon93vSqGPxiMNG8qi6O3hz24uE9U/T/0tv
3EWDSlBLkCVrmcPjVpcj0P0ReP1mAbmyO8M6Zc3yaNtoAmyHjbO0Tct01o6j5XRcuEXSfRm+gxIR
6jm5pYZcXB5EX0d3UZ5mGJegAPxyRnLrAjpYApLjho5NUedqBODN2dAdcJO9pQLqfOmv0osjb9h1
7zXwgq0K8kzTlPEcETDb1CFhdJVgRn3Qv7imxoKFprHXUxRaolEMzJ0+NNLhO/zxv6KR/pMN+8ex
fNeqHNCSrHJzOhuXJ7fhMxcnJtmGJOuMGfbX/A1V93yfxwyWh6XhhD9xPowPZVTz9K+7L47QagMb
EKO4cMyMDKnyjbmZZ5UoEFUlsmkQhB2dRzjhzktKHy3+Nd111Ymyy7kfaXnROH4jwlcm2wXeVQ9O
q1omu0BsAFvB6osSjWWwblS2giCCZOXYT+LyaWxncpszop3nrJPzGe6cvtOagd4ShPwQDCgz1sWP
hBYSFDdyGvyeQOexK+CJHr10fjlRu72BmTbffBgF8nBaRVQVBGyE7doe5qZvbpZJRJSb7S7z6l9O
p5jdEnOaDPoy0R0cgvHNtQI9PkNxrnoKAqIx2wR3OVZNTicB2cIn4biThlGAqkXkMqepYwZ5Ch+m
XE5knq9Zrk7lQR5aq9QccQ6+hwg/rRxpzWN8r7s4IY8s0qPR4Kg0g5lzPIAO7zTsv7nyzrgxco3a
LWIkNW/0jFzxgFvnLraXgPUrATDrzaOB6yJTSnGzAotusnhSuJdmNlsfFV/yWVm/I0zs3DSEulwP
p60M8FekbFbjovnH5HOqHG4NjvHHAw2bvSWOYiRaNm3Daikj7+LyZetuATZ//YC3LYmGdHlPwykd
N96HmcZZB2abwmJQiyf8MqgC37mKA4Psj1RR1UBXFhrdA0/f5Yrk6cX5/HTR4o0OR6/TE8a7oYft
U2/gWD4z+Wr4r9h7yC87zqJ2lZftPlcsHWXgn5HCq8xc88UJzSTEfUAFUy+pcs4S0AD40oYQzbsi
5n5WKlHK4nEEkL7N6dHyk5KFkunHzqu8CrwmGqR8Door0MVWBwIH3UoFCNtTfE4gbuELspK5D0k1
zuumqqKBvuECtEamBf1kwQn4UqmpC4W0tcfG5wMjU5oQZAUNkAyDUS9cbzT9PrX9ARbYftV7rEuT
Nv/2BXFDCVV80mvfz7CPI/9EXkxJ/VtX64/Whvx0Nh1+hhw2OJbPRd7KYAo36+8A1DUXsS4h4xtc
/8Qi2uaiysPXbUMdSzxRNHPNrcOp9dwXeKUhUdBIktzjRCAyKanwKGos/V4eYXJxbx9u4r3vJ+nt
z6r43AaxnclwNi4ly+PbrNSzCd355f6OCKJNHJdI9V0e81sj53td+2ejktXOagLdv6rTsmJpISwU
ojK1trAySbRv5tAusNc0352lyW3CPE/0Jy7h/cYm3La4DzMNvfv0RrfQbiBTNA9pVJGlG9EEfZwR
nK5nf6494Oe0+mh7dlOZWzZWdl5jlJuX6rKVH97M+4A48GRwfcCE/g8aFrKf8IH7rsDRnjVVZZDI
VcIxsDnyaBh2BWcIHGQnFLJptSFCbFhOQb+UhA3BXSVkWrMX2TQXCLcavalqvSsascjquhBDBJV/
5iSUsyiZrZLurWsL1+xONKKf3/83q/tua8rxIvbOkqe8tlVS504V1+mOfqDFyVrRKc5148nekBUC
Hgktl1S2izBmjJZHNiCB05Ef9od+hMabVcNVEIDwZVI4EhbbhDLD4gTk3qRVV8AMf0QUFr6p25wM
dmFW4b2Eo2cm96AzckEP2xvPVirSO6WTVKxEipBzWCTF40HMplfOIlZktD4fXvXG4axFC59NFh7m
wlBT99uWzyY4zUApnP6+1GQnAmNyC372ZhE/VvShdbnaqByVO/OUzsGCOK5+gLitQhh3NK6VPdKL
SAGQpnkhiE/pvwHjS/gjqDdBOnTJbk68uZhu0j4sE23UwFOOhu9mTadP8ExE1o/BdeJkDuDXjkeW
wlPpVCHXp0E+mEtZazUMjHHfUPzA7VQH7m3R5OtDIhYxYnklkDqA7XRxXX3cH8Y3NW2o4K3WHVsr
wNDmu4pObdB0IHkqsPzFRCtNmG/FTeOzyQ6pQkzKDwdU078EPP6n9GXDiGZtkloTuQLsMxOdVGfY
t+U60ALjpbCbrgQilOCrZouOOmRtmzqqK79De1wNSjTwwwHeJgF+b9YpKUljTiLMJ/rPavk5Paqi
T0XY+3eQsfxOwYaMDNZqT8WchVbX3FuKdZM6gE0r5nt5o0RjQKy5ALFQCzttbwTcmZylBOkGsT8/
/tCKlsV8VosnFc6UKheo7R9P5Woki3zL8eQmebmIGunZLTuiybvZ5BmMk8+PxZJ/b6lHj3pNO0pP
NqJ/iaT58lILuwobGG33ab4IdlMgGCSVsy9oTbxkGoGTo4KPmfwT/78yg6LDIDzxNkP32kQNiOLG
sPbwhU6wGhwGc6hGEJHMYjmrAEzDaer/6ryY4XUubf4d70fpf4x3n1A4zRpZmnSO6cAiB7uoJ4FY
x+pY4Z9x2JWRX85MNI2ZhzHtG8vPm7suVySwsIwqn7yv+JPKtQ0xD7Ad9MAJveDDj8f3FfwHqsp7
HEdYyiig3QAeXvOgplq/3VjUk3W8HO5VDQ7ASpOnFhnYRCJ16f9UuH3fYWilZKARjmguU3TOJx64
PHarKz4ETEQU51gwuRh/jyzMzC4nQWcWCvOCLtQ85D65uoK8vQUsHjJTzS+5bmDwWfaUVARxa8Sm
/VzxuQohzLi8NKlPxM5BV5FP5iVOYNtiPCNGTNPpDS74T48e3l/z/SmUhJDWXHK9gJMsSMmNzY7y
D8PbfSr/mYuTkWkD2lDTyCCNR9EWOTPLf4GPVCTQDcp7ZyynANhHCMpTEkOdN/08x/qln6GTFIQ/
NG3AqtDjFzGnQSh+4BEjheFjvn+A3+i3VKhR7V6ZJxYq0p52dg90OoPCECwd1SDn4r9hFmb7i2+o
hQF8F0YsLsqbpFF+sUsNy+nWkituZnmgTlB9lbRc2slsbBhBKhQXPGoq1pJoO4chc19xzcoBGoWw
yURT8HHIIY0DxEuI3AzLukicESZRe72A7lJpUipZYTHgEt3KbRDbzXm2SSKns0b4iuH+jUTyptgj
J2IgYt25PbsbMRHwwFwx639ODE4vrcRy17pObz2p+2/mLGk1ZaOHYJ3mdXxpIbaFnTk7sLvsU1jc
fN8dQdzIUbLXywhBOpBQah/NQze7hRbEHDfKJgcRmzL83SJKe0Hv8Yt71W+Qa7sKFyZgxPbRxE3W
EjScapFOfu2BBM96somI3WffyDqQYKjPDc+0ZYlxAeKX3Y6RsxgWtWo+N7Go2pGUa+9vrktn+5KL
0xHvqVXOuzwNJzspRiDbuo5m0yUDinuwNXx6RyUycjfvUYve62ILhzdy8acb4uB3KHsvOA2/bT7x
tI4D5apW+0bQT2X8Ah/VHDkV0CliHx5+1939XaLvAwTstNlFAyw7fSI+MfnZNY+2aTOwsTlO6/+x
Qu2odmgur98YTw9FjN3vJ3uJmm+VBwqFZx+xSmXG48DLlkPbsw/YpfHtCBXCg4f7tw1qmavrVgDK
upHqj7tb8JdsOPz64qSvtAI8GRzKppZMnyiGNxHKb6uI7FPZjOBaH/ohSIafsAomO1AuLA3yGPr8
Hdj9fm3ezIHPwiDM3+Zvs3WG8erCGfvpyZ5dZQuHBe2BLpYiaWwyIY590maYtqwSIT6p3050A/vL
85hQQ6NZ7bZazII/BAIN6Lk0menTsycQdzjQQiq4jZn/z8SwX8ozadbKZY28k83wp5sN2iS4R+2j
5Ojbp3YkN2oTO9TPOgAqWs8eIaYzwmqAd8LQPA7xyAEd19RNIryGfQ6xmjoLB/Ygbppy7DM6mbh+
NKjRGBXc2b+LSowC0jKGv5ElpkgmU+IYfTIhHb99jXSjOxoZt3xSW8NK9d6nQk3wsyw8lO6p24sE
LUS7qqtw9eyccVae+7+Eq25z3BqtmLekcWM5ohp6A5EBecr3kShVUUy+vFvc4mstAnm34EIjgS8l
enTm5PAgXR6IqmFwixVYETrYKrXOGakqqxjTddZ2Ur6ZgZ7xs6So2yD4v3QfL4iLD9bIOsgQaqzp
4uHg/d0qSjyNKVTiinold33ezEvS1tDt2+Xs61+TA/xw28Y+isNLGOkz2n7qEKoVzKvtWUMOxDyi
C40CXu9Sqafr+3FB+x+ccaGcQFqkZDWfadWEcOECVhI/KroLVPT77ok6pqTY2hVae/ga2x9+hKdn
BjzNsalEriVGzpOkvZCiz3Ry3k2izxW9r55ZEy99myBKIcsg4SMCw4Fmc4KsrFnB9JJ+eqOw/Y4s
D2xgZooYbjXlIkOq0RFPlvMUTbAgTb9TVsv3C/vJ+xQSWSip3uSXqCBqJE9HaFipHN7B0Z+N6RPh
KNmICgUJYVRPjYtvdnSLW5ZEnXXdJUrsmL4alp4Zq268t3Gly/6LmpxPhA5qCICAdl69TfkIMlYG
3zscXNS2onT1Ex9lv/tFyZpKkFJLl+z6QsmLe0j7UsCSy2m5xeFdTd/LVFp083DKtMWgA0KUErjK
WHAeToAdjTRkf3HyTBdI/fmU9ZTqf9GU4Pp61ql4DelYolPdF7CGGYvvt4phBnl3sFBdhS0ZmbD1
4Rzrlp0SIRfkWVOQyS7r8CxdJCTew+c3TwDd9gdN2cMTiONj0hAuK8p2RNsAHGf1vvxmaJeLWhRa
iRSwjaN5zTWT3vG6976hGoElgnoKLDPsDE+cc65h+ZF9p550fSEs4hSjfG3esoajFCA/pnqR23Y1
44iAhB0pctApdu2/4SDF5aHJ/YcUrKzEhhRZXNcLdcYJa6KLWCfwWcxcINV1qOX3Xh3m57PlYQnJ
qCvxwnavl87SZRkz3NMD/po97awB6+I92FmUadPRwBRegFRMP5PLUqyfyYOeYu+wuc9E6EaSv/AP
CsBUAWkEJYdZQvjI3oymy82W56BhiY0VAAfIw4YEunPr0u29sawhumKJKFhZW1f1KEcGhNs38Vsb
re+jv5ot/v6c93SDIWD+CMLtcNte7EEW7f8rYy4BodiEPHbopZkuk0MgYr+15nwtSD4JJRDtcr3O
zqiScviWKiA/JIGx5DVctZ9IVzThFXlQ7RgTd9Gux8z1mCTVG5D5skSnK9YW7vaHwJLXTkgPL8YR
6sdCnl8ZxlePLvp24XaaMu4igL4M1O0v3VmYbzt4YjPhl/FYOnoYiUylmF8IC1KaFQgfM6Hm+2LR
vSfRFHiqJhC4jVflRnVKztynVjuJg8WFfnvW2s2LK6OmM+ZlqwOcoMpqgeeeqe0ZmVzhvt5H5BCE
FG3BTx+1gCMCijTFLArc7dMIyBKQf7TcZPQ/ft4eEXSANhk04L8Apqh6FsAuGV2kUKkwKdOr3VQ0
hrVqbYz6DvAsxpfxgvEkrEeYFHeStnCrpRgmEliuytcLpKJGFsN6eVK9b03KJGNI4NZpOlIfhWk5
O7oGmjLvrYnFMRCuOLN9D8ubcktoCb5WBSHtfIvHEHj4akOCUqd3e9JRx44lPmjuOO1GrBAP/Zr9
N/nYgyd9JVXnsXgmD1S4sewZHk1uxmVSbxX3mBQ5oa60Wu/fZwJ82MEigjlNspO3EPBDVQFLnAZl
A7+zJfZJ8qzKGh5MIq2aH4JE0FtzjcRakarzwnu5D5WWBWSZdAG14NApNBjphKLEEgsKb3rkPHIq
ibjHOJdzDS+s5+NhC1BurvCmRHX651CZ/Lp4c0CfP4yZMuOL2I+MS/5rXc3C5NJuo2F+NF/bLlL9
4LzTUZRioOu6VljlIjfB4/Nmyl2fuykyDuBDGesTXw+xQt8LcbiBUTMArPHkL+j0lULcnTOX0bmK
RdavLXYPQNZ0iMXrk53c4h8FUhfdfhkeffmggFfHzeP9ZNQk0+TcwdKTQx/xWWc8a2WToJ6lvrw+
uH4yF2XWqyN+oi3TIHroAJw1ZhDUNHSSa8qUUlXmZt5I0HdGQtPrpnHnUenx7v0WgxDgjB9Hg6O1
iVJHepVPOD4+rHtryITa5EJRtJzsxCtg+M8WHmPczv2+z+G4rnlvvdkFQ0NxkCvA8akaryQypRfL
dma+LK6YqmC7Cl3Ob48apq+H0b1bOAXNyzR2J5IvXT3Z2HCIBb5z4QGm2B4mP5/RYNBrdoALcbEm
2hH16NxWmpATegjYzU5l/vU1mvgq3a8KnWp1CR7+qsekAD+x0s9gtt0liFLRjXl4nM+ly9rgVTTR
k0w1CZJX1eVAjYXhlGZOJYWohAXZAbb+im4aiOEtHzJCSr6Cb4oEc7Qo/igQ2QOEVV+ivMmR1UQW
zltnvoglFoDEN3glUUguQKTS5enWCYHsAMhGpdAlM+8mGUXUH68epAxHAO9Dv1CWJ0mhZ6ASpCuJ
BnMcDcD1cBqMnwJFOAj2ONoGCA2Ie7D47wkJ88Lr9/3n5OesLcjyrd3HjfaTdFibF3+y1tkovLBh
dvpS1Z+/DSnt8Ps1TkvE05J//N+682RNE+zIp7e7gO0qxyCQzqQYcOm+lgzIvw0mAV14c+Q10NnO
mSoT0paqNyaLx4bGnhyEaZkUwIjSGr4x0RGXOn6EXAX+co76MFYjfc92KWBubM1EjXD6EtlhQNjD
vGCer3rJJ119n7AHW4SmpNbEcYWIMHbyQdOhuI+y0uvdQpnzvjOsetqSJpaZykM377rwwWJA6557
B3Yx8jUkoafuJxh9m7E38JcN6J4ieFZzu4QmVLHYwhnV1fj4AxBo3wJAQs3PsEcVQXDbCIobSaT3
xJXr7eL5lJanF46njnlDgd2icnRSMj9+77Y7kCEyyvuHkmD3PHHBREMy7ve/zaSJSmQAQjCk/YFQ
gKe2ZbkJfi0iVrxjfHeAK0y0dDHCN2K8SQnh/4PA/RkCRTj5FdmBbcJnHv98MGP4zhNBwH2m1qsX
qnJoBsdYzIUtsu7jn/UqFss4WyYT48af97Q6njT6w1qfeO7pF2KBztpkPrCnEDDYlr6BOZl0E951
cjZxpE4p2M7gjmKbBhvTCn5E1fFM36l6wPPNaVRmGUmsKUCmyZvtlTNAszYxDLba8P69gz60pQeK
q1rmNUHVIDsV66dstESIr8UPEryU1H1Oi8Tap9vZc0zZv3ZiSflvUbZuAoj+5gUycVKOn/IZeOFH
XGFTkPzbXsJAod72sQLQsl0P2UQAJHUFeuZSpIN2jnusBZxix/7tUC7hw6zn/GfzcXBo8Z2wkbdW
WQu1g1Bj5EpT7X+OscIrb8+dVvwrt1dUyhWyxAxnMR5laQjxlk/4hwjihi+WHrFxynqFtxds9DMG
vErQP2P0ruazrc8oourV1HFUbe0/J+OzbVo7eqnSTVYsJkOX6oITzCoTAxyeXTBMLLlmQrmL/fYt
e3CyNqEArXIh/0mi2j3NDDiqwlfymfEDIxJZ548/kPtsgr418Wy/nrgvdXW+00JQuqgY5KTV9dWf
7uBpN8/8TtHnhewhHJXWY9Z77VAiki/c12jabZ7rypOVBgZGHv0+5HHT4NaMpwMg5IDeeSxskzkJ
ppHKYPSizUgzLZ8jAkgJ48sCkEWnJvPHGzAbgjF5KnzesU0uYa/CG1W7lSkOYB63KBSaRR6CAyoA
AKG8zR5q33e9M7PIDjoQpaJvhtmquOyxn9EVQLGPg13IGMtZj0ga4F6eEQelBIQE92QfjTNVQv4x
q9pPNC2B7cmVf5Ede9vJEEyCPXLbq7Px6AhJsNKor48vytqg+I+RhjX9YaBomQSFERRrst5vFm4G
2jGUXd5XFXBZuWm56/VL61JHfP4sehvASnFU7DGESNfIhYNF46sq0hU567shEGaGzw5zZxwdtq49
xIju6KTMt/lgIgReYcwXEZm5er8WdJ0lxBctGgjejRBKHqVIE9odZ85Ivgxh9qFm47Ejq1iyn+6j
TqnE7ya7mdq26rIPlebG0UCebmb2yyrbB3xNpnci+nBniStGwNWglwW2jBum6H2ZfpDU6kHwMHDp
Xlz98MPfoqyFnWe56oJzH0u3O0ys7Ot+2T5j/T0xHhBvwUbFCAfrxU4Yr+QmqkeOKrCJnUju/H4V
FeeM33C3rKzxWqWXPJxAt8JUaH2zntmCuvBVzaT8GyKT3IEFoExtGwe2OH2dOz+40YS8w7QzEnAl
Ac7Qt9mwgiOS6HvwQ5Rh0IiJ60Ha3dy6zEFtVuIBK/tA+QQScm8l3GdneKazUwFSe08CRo8vT0/g
nUMao56MU7QvJysYcdAOp0aqH7EPgDFJZMVSjIORLVXVIoSZD+ZA2r2NnO73+D5/p1L3mbcitIG+
CtDctLkkIGxAD9cuh7P81U82AtS8Ltk/kw9/0850ndvvt7OSLPE/IQr5ZWlkv8OzdSlRePzQQROy
VBa2efPvNJhrws9PtFUi2FcnGwyhwcjAaRyHC/oCQhg4ibbGOMmUw5OK4RJAMmY/14mYXcHvZ94U
nYzY6/9KCxQWD56S8Cup11gfTDlQ7gXVZZdMzhiHY5yrH4x1gtxYPt+1k07lm2sq/2iHd9qf2hy6
3DQDV4te6KfI3PVx110qE3ruFclDMkPIEVaunaLkuh2CVrDY4IYj9mtEFYNrzgbgSP6ILngpUIX3
Z8q895YH1ZXldGiM5VyxkSER93wDbPo4+vyLb43OGG6Bis8pZ9Jrn0GcKIF5lIgVqso+p0il/cSl
fFyKx4WJh1dqttTV4OK7yPqpWW3bc8BI8LkG3AYDpeuJ0Z23/MLYJVmyLpvfLd9LAlEKOnzKqbyU
+40muJ7faoBclj6x7eDiomz4RgM31Bl917Gt//W8/3FEbULFnIe1LfAL7nkudXevRmhpZiZ6YVtk
8GlBBYPMQQt6JyfpZwjxZp2EpLg+3ZcRticzb4SBdJczGRJq0xFhoNz9TL4hJ6dZbQ6Am9fIZ5FC
Av9Mta4D7/Xt4iODsJld4GAoe0JjHsmloaZX+chhufnifU+QWjilh6pl0yLA1ahgb2cdti8uubbv
9U4fyuga+TtcKcxnT1Yutz0fROZzJYGk2m/RHxIiEffsvcO4SMadL9rtLWQrjTS8nHgEx2uYJJkS
x7wkQyl0QTPjebpuudTqEhm2AjkD8f4vGnNzPzrlDVIBbNtGK9D4w4JnUB9Vq2oXDTjf92B3VMUM
36kFvLb6BZfC8GsqZn+sQpXS5xumc+UO0OykCiXGk455z27jaAyYE5n4C4d+fa3txMBUVLX5B/3b
Rf5rqfxZTnUlNXBjYbWMKSNSMNRJ5o9AKcVU2CtUS+3W9BzsMrmzhJOm3Z/SZJyIMBop/7zIyk1L
L9Uvfi1hOvY7NZy11mtVRsuieQWARZqcAeqhpMz81wGpCnl4WOEntBqWuLsfT3KSQe5nAxBJePr2
J6WqXQ+lmLC8IJ7UnoMFNKPd7LxQvvgQtCQSZs/vetOH9s6Rgevf3dSvUQrqpSiw9mWPY+MyVrlt
6Rxt8YAUULI9Yn+zHmFvCtvmoJN1QWKs1DkCSdIblbOdE4IemGyMBx2ioBPBlkoz4C5vpKvMzPp0
MB6rVdhvapcGdiIORLBtDclkX5jxh5x89FPvnD6pWd0ar1xaRYt2/ekGR6NEpi9a0cepp4jo7Z2n
d+U82SWAHYbRX9MnMy7erkfWTv4mapP1cCULTG791Ck1B9Ew6eIkLOaZHExVk00IuwqS8f7hK06t
jVp6MQR7P8SR5+lE9c7MSaWgdhLjO/M3ZP6TRdqD01+Gwg7ZlsGhfwp3J7WaiCEcwjtv5OBHXWni
6SCdrwUh3GY4lOhJwQBDN8CHfZKS3z5ZyBpjyoZ9bvxCjZQG7ANQPz48muaQ5nZplB58RcoS82CD
HnBf4TL002pfCXUWFHKuPPMR4E5r4qbkz6JQacoytjIY5eyyBN51iZ1o1t5a5aQ//c0FK4fr2uNa
VxMLzeqo4CKSvOk0pwZX14d/VSVQieOLcjequRGEcRvJczijgsed7ZoWzwkIbVAf3crkv70zrVN5
MneRZSJdVozylWeG3iiUHZbPVCLnysRFqjXEakvBel4nFGZ/pNg8h3Dd4cCNPd3kj4vjQmhyXdOg
5TKuL3MUEdtFSv9nWavrII0GJOFWl1xTXhfuI9Rk1H+ruVLY5PtyJWARaRKE9X5IxakwvlsG69ZE
e9DPHOHnTk6f3IKPZHgtCLBpwj5ngmnRiskzpY0n1cIelvT/+E96VM+FTcLuQkwuLIgFGI4og7EE
nMqVP4pS5yAxzG8gjIs+XhF0lgWFZks0JWM/cgaDuVl0YT6fKtM/4tRQsaiSDG6oRhT3MV6xx8wD
sTiK6X3E3oUXmdv5/A0y5PB48KIiGSHf8nVWw3NNpZHLC+7QSTn6HZT1qiIn1oUx+0qX3pm4EGnN
/0uOWSQJB3JeGRifJugs9JDNqpWcuO6TUZC3ImzKdUlkRwYoh9uLp6qeGSAdsAOK8JwFxcOdgkQb
mKlrkd8pBazXDxhuapCVq1xm8FO+inA1TqZbXGEGJl0TOEQ0nzei0VTUN8SG/0n4dpY/tTc0jUf2
z0NLrghw/TJlLE54U2slzTjtsmbGnux9Fm8uVcT3TDjI3GRoBCdc/WQ8f/AV8A1i0GMLG0ipVwdM
2xFrRxixXiJg19gcrrAgr1Dn3Zik4gz+Hdb/W3PIWZ5wK1l1VadOnCSv8tMo2HpHG+lNv5e3O8Ux
dDVKuClZ3VVVrGAnbREEO8pfZDa5cIPwq4FhA8XkxWNqzX3qMbZl7ifFyrKsi/Jwtk/Pzson5rO/
JoGpytFCUUevKund//DCalZ6zOSOgs9Psa3b8drcqKJ5FgMnYYJwrpt0DH9nu5zXIxwJG7qN8JOp
+P9Vzhf0KS62+p0EPjg1sdi6xO8HibwIs3JXYC0wdzWGsAN9mHo+NZcOzMa742MiwIwLmy75z7w9
Tjw1mVhuN3em0goAaNopyhq52pB5Dwi7ivzm564CNF5gZi3JMz31onZrtbIrA/fNZcw6QKt4Mzep
XtllhE5MCVS6GpMq0FBfAg97R07Rqda1Mwd1EK2Pi301u4vkZwGNYOIUsqwMPrEOo9X6jowlydZT
oxFYophSeUBQPd3plRgEi4D77Ldp/nYDke9hIicEe5QIZEeITt/p23sOfUIljxYTydRcy2VZLOeF
iiz5Xt3XRb2lTgYzRFErW0vAXsE0UJmuaD6tSwSiTb2Sa2Bjavi0IrxEP3YHk7/z2iauhyW/vSEM
Ip0YdsoAzC3RavcWiBIjpyLE5TENKalvw9sow/Ah8mVfdiJwJl1F9BgAgRkhIUfKcN2aOBf9x5pU
xL/iyltmdXc6KfT86OL5lTZAZqdRNkh6CbHO7MiKEPjsBIz/v3Dd4vIj1N/0XamLQgOk6UdyhiYU
+zGLEHYEIPmAlWWc8Tz2y8YJbeIKTPeA9GTXm7zdz6pZvFrLDX/9ExAv/yywnfkPVbjoOtCXoMrV
6HzmaYMdc5rBprjtHyVZAVvum5/fPZZs668Qzy7pp/nNnpwA8ci0cuESuCF9HjE86hkdD2gZ6xCV
S+E5Unm9St5F/L2bPvl3HHvFfqNKjnSW/6zzJoOpXBO35kTpdH3wRR0NS35VQccvCFRcLlT8tUGm
vw02/4g0QcVVWiYNXqcbFc6MlXeU6g40Y+DMWoq+H+h2w+pJzakV9HXoaLUOs13IvOlyRaUir56n
Ys4CX6kien47LgIueWUUh17R2FHFouczJBARo9PZAWZnrBTW2DMSZd1zG3iIbaRiSmYJQ1sWsK30
h0Qa2A6Z3fBuka3GJdw9wDgENb4RVzK1qhNWfECIXWlCclGWewblYYsg5g1kopmDwHf15OD/vODL
cn2cU7wpQdLITNmSRmm8HQGTXRJXdA37XUGkKct7UW9KLXr6ZwGLZGhii6YMh9x0zEpws+iEQiNi
AHOb7yD4LRnlDQNNDqTYOt9RrgZPDx3D86iStelabo9Iln8NQdLr3aB+b0Ze+y+2+sK7AuwS2+q1
Gi7o6eSfF9PKBpNdzT53vHdxHlkG512nTPNrMwMfxDwFJZ0edAnJoA8yuYR1sR1331OAXzGah3Gj
CoJPbhb1rH0rXUiuCAgXHi8ajbt8ZPJ8gN+2qyP4hPLahEabrmFKNP9G/A5jwJWIeS+FvexaGfie
NZ+mrPszOlv2IdlVLmmVk4+UKdZFPg36wFXV2uSNcJ28BtWDss5NJJO3wnZfdZ5vZ7d8246xUc1h
0kTPG4zXKza5Xd3JYy40LrzA7RV9hGiDsS7/oMkhLP2WElFWNKB4WeZSc6QJna2ltFs49Z1xb9My
VhMC/e2SiIVjR+2Lgn5WJOwJdRtTEZToB8iNjCptuQvCcU+fKcZWDBhNpRp+VUPz4eahgy7I3Ngz
5jVujUhve+QK7Eh+7Rc3VPttPu3/QhzPeTuKXyx4JNtIvjKrLIGQUJWg2xMTSEwpWPJSwQ+iIKKa
NEzYIQKT8C+9+I9oAzKLoSUkThJVqDNO0u8eq4koD/uX6T/XeCKqVacMxX5y+qnDuFRZOBzWpM6g
VPnGHAs7jdKv4x3R2+UMyBho6Qr7o8lNkFiwOyQzquziH+Mbb8CI4Xt7Be4kmRgdPLKMWpBtP6hg
XBw0YMltyoAhqNBPC+hMCmmcPBczvE7dsvLkSXpwAFYreAumGsJggsBhZlL7kXS82qs+EhY1V42P
Yf7bSgC6/200M9wrG9Uit+pYbtW24VKMWxz1fChnO+W3r+7jOTGG1C1QW7Sj5BDhEEZWx7BGAY+r
TrKS/QqdrEoxCPWAmTifH9t2ukT8+P6nzu06FKD26/sqFcniBmTbOund4KXOSlk7bcGComJlFf6I
LVq5IIqq6TN9t4589Tj8b4o8wzL8tc9K9lfnqYZDZwrDw4+dKOAwRsuyuGAVc6mKAu0FuBNRtIGy
+tj9qY6C8sgEjlf7tIs0Hx299IdzrFgzw1aUe9SYoIfCcD2GP+R481kPkKojHv2k+dgDMhqe3gBV
hmlm0cOpD1WFgZdC133ZNruTUqHE8n+pCWiqLstYmLDIe1M0ptHRwmVhHFTQ0nqZcWav8GwhGYVW
IMXkrBKOkCTaLvtY2wUtScPigIrmI1jQfHQr+wu2fIaKTkJ1YPIX0m4KtBiY2JXRTltDQWUYdoC7
f4VEkcYIBxXT2XVlycN7fmP3d8bjH2hHfKHxCrzfxPUhB03hOdYBF8/GYnaqChIq3YK9QZiceN16
m64BYhg8ZZ8fr9OxoyjkGc4MSXG4XEk4WH9yADDCEiKK+fefsriskoH/xB6snpRwDPMOvnrBPOme
I9jXzImVNJZ+WbLVcWkSQtAh0wrtK44oHzwtx1Jf3FlxC2B2juBelO3NRHBc37PF0c1WHC9VgXic
+BUnfO4HuKZhZlR5GOWTSaWGZzBcaa6f+z/5tV59WsBYbmoA21mQbK6XYkl+v2ZAUm5QEX+gAhrx
/ZcvTHlxESzmL4cEOpJAg9VsDwrE/aCHJb8V7PwXxr0UHBZj/BqxzL+ENvmrJUf01S82cU1uEQyk
dLGPdzSiCnsoU9XFfAyYFN5ydq4UbhU5asa01KoBXYHOcXJkL5kQ+bRxdcjTUOR9Amn2pZChc1ui
KVH+9UZQDkZBl3kYlDLhbJ8oYZYvnCeQTBiyo9TzlTiUeJXEWznReyNviZC7RqEyCbFgDcKo3xmu
ChvMxm3dTof1lXhtgU1paJC/6CPLQ75suiHS5yiVIMVafpipdYRpRdAop0R9ewUTNfI9i5h17Iuf
3XaJiLk8q0srtnaJ8Tbcr/8t9MnpZthsusd2MqdPU920qMnXCLkvrhUeejHHEVpiRlfiNkwFHmza
LKb3nqkn+BVTrN88+qm62Hpd6RApXVD7/tHi+Nv4ZuaFtbUgnhTZMbCKGas6un3VcEovzc305HkA
5EKVVK1QURlSj7Ab5HtXCBEJ0msBSSHnDwd2BIIeBZtMT5mHiI6ThgjVhY0ZiFlVziZG/iXAB550
X+XvMLo5bJAUNaczyzgOZTRtWTQIOeXvbxZyIrFh4dCYGv2L5h5JCG6Q4wIx1lRVw4Kirvl5SXx8
Dxj8st96T48obxfynK7leFIKmRkvdP/RfFE08OGk88wXtNARLB2046lSkS/vN76DTcPJseUHAQVq
Ovz+JTlm8L9O+aVRW1oNWfVTLwAumq/aRRuUv/hStpn2TSCWVv4czWscafu+Eq64u11Q6+G4RmD+
VttLv4bQFOesyn2Dy94VXE7DtbWioPw8MKiQjrC1YBeoRZuCHyAwIv6rOgoi/rP9BMm2yYH7cQOE
Kuv7Ywc4uOyFcITHhJGTzqnJvaPRIYih27tUGaH7EogqqaTOT5H7YxFqYYM7hVsxcgxk7qXxbJYN
EZ3ducnVDMQAzGyYBDUY28K2MaiLQekex7GGir4fqS2HkZ90nTcNUJfaaDwIAY7IQLbfVEXIfFS0
WeVw7mb6QE2sY4bYTKw+6hK+6q2zfanrw0ML//irXTLpnFzfy8b+XkwviTZ1AUZkyyjSa0UXGNDh
d2iOm13LH81DLqMAWoa6lC33L0sQkSK7vRWsbMz7/okXgugNzp7ggx0iyrupf0/+afI3m1vHYvAQ
twVAqig0xD32XUfjVfY8RV34sE41pDeURD1gkbZoHLJCRQmjui/Y0QZlNUD1DgnHiQcIstbzHHF5
Eqmn2fba9YQjA4xNb4quctQobM0HoarvOe8+VJSvxjjugib/ZBD36rzRdootiLnY897MXHNmbLDx
EBxGmRgr5MsORxum1AhRY02RogC4l26OUi3TXeKvWaDlgEwOUwg02nWlaZNWC6XPnZmdlWBZ7h8m
ilBTIs0w6GsPeJuls3tKZxmS34cVherNCz9xC/a34DTwvAQffVNrT+VyYFupk8db5ZKZQOlW/ey7
qNH5aZ/zWR0tN/OGksDFqAEWDqfb3CcJYC4S5mFg8ZGuJuksJHi0MO+68TLfDWjAWNhbLBrudaai
uZ97yl0B3BBssGOC4Nf8w9lwKsWYevUhNM7pSpQOC8A28uYTY44YBpr9xI9WbJEYBdUwumjNn0sW
ykUJ0YD3c5KySaT9xt53bbnMUxEdTWmj6VHE95xPmpHtvo9E1qxWs98zRlUirSqdIENQHLkN5UcJ
KZ0/wX1wrKtKrZYtFaQU9BPH/z/NyTBoh1eIWmAH4XB88dMquK/L3REHzLHRNVocabAvbaSV3pk0
tvBZ+gn7yaNAwe4yR0aDcQ+8NgmPBUVH+skcDo3J+NDHonmh5sSPCq6aKUCg7fIKpN74Sy7bzyJH
wf6yRkGchZIrL/szamdANgv7mx0P/JJNc+4D+EWmp5SlEKrtES8XLbkIP7VfFdgKd9sfj4L725SW
i38uhg8X1P/rhxWnhI+0hbk7p8/DgcJUgDvP0RMCDlG10pFp/hnG0MZ2J6oTaOD6QnmG4HWPoDgt
7bFyxUknudz/69QQPTITyjDm++KX3F76W649PQBCIdCjKFsgIsJg6DFWlzIiLJlr3ePolLkaThx/
0rf4vPmPi/Kqabp8efp9+J9OltjfaAHWK8x1FFoO4nuxBlgR7Q6W0Q5xjy7Kd9WAHcxFN7UUwBdX
YAzNMmKHEy3JUbSShZoYQKynQmh1hcJYXYsKxLPQWvpUnald5kK61MmhmrISf2boDlN6gizrxk9l
1qUVJ5cgXcjAD6qd4WRN0lAF1V6uzIxhuoGEgsBamQy/OolMYaEe5vJHpoTI9YMWARFXndVT8KVS
7qpbRYC+1zb9kZ1XesmcTY6GlApbX5ByoKHs6Pr9bsDEk9WxXdUSCd6C0AgSgf5Qivgks8rI3hFw
Jli1/OBbPjiUcCohKlejCJIPrs27NDDXeeIM8bUfXRKeFmLd6HSVqSiijbx2Fr5eD1ywWT8t2Hnz
XkhYq1toLi2rlglF+FmOCXMY9qJZOQbK+0pSAqrUarcqL4zPCAtwsMHP4oNBH2nFVZuONf9+j2Dw
y5LDHsrfLhoLUIc9LMC1bc6dzcSzzprcnZl4l8EucFbo/Gx14XBnRpMRRkTZ/d+gAc3/NQTTlZed
w3HYb1YF+q5y1M5VZQ/I7Up4sJ94ZSPlfTg7VYkw6AQYEGNdo73lBGSoWlD885r2pnkcnb/FHW69
DvpgPehypHg7R7xbAp5XVUpbsnYeW+7UKQB6juoV1fVnc4l7Nfjih8g8VddyY+IyTHlOizUYEIHn
K8Pw1UFnGym06hH9RmZqdnokxLG2vRML9j9Eq7xcTMEJDyUbMdWkps4FyMgKGy91Vu1yhOiD59fg
RG5sLGs+6HvGye0qrDo0EYLXuhYRHs8SYCHVYXwXWW9QvvzGXe7ywl/YSvbnw3N4OW13zsu4R8uL
Epfz3ed+LVaef9wyWoWMlWXNV8m74uZKcTuTRV4+4N8V2EAacuEsyxv/zV9Hw5zlv8ZYbNh11mbH
XG9TTPDv2AqpmTbdwE2iscNIc8nl08QAiGMIPLo8PGg5RCXHjf324nKNLUW3dscDMYr+oFSnMUpH
9XuGdqQHjfxWgo7sCOueGj6ejKILT/jqKzbKJ6zXlC537AE3nmuEPU3HJ6ArLLVGRr7H5R85inuN
qHlsC92U9KOFZX6rykZ58EkRvQSD41IO1zNFx105EGV7KnRCn22repKiacRsRPCuNIFpSJDvRYLP
DUXcRRVNjY6GiNpCZ79f2Lz/axERyi4SMdUaCmzznSemQIwJ7qiIOInaFqUQ5KE6tzgE7xpxRTsn
uWRuiJn2YWM07mEAk+We0qyizd96Ds3FKz7m4Kcl1vCHHsVNCznyy/+7hLp5eBAbiZHIcJ8y8ZQ9
AUkhKd0JgRFDSvCaXgUN/twZdRhb/R7Fa4tfV5hkKZL9UnrtP0SP9PdeAsdbczmBWeCxudxNnb6o
uOPNzp01zGSme6zuLo5pCmcg8Rj0TI1ubdnvpPmRXvlhe32t3V0pnz5yC+DejqydrQGecK6UIug8
Cv/FkrB0eTJ/mawie0cXjoFt62O0Ifo3DmRnCKWRiWj+wkiqpdYNurNHvgyIobmobB1+G9Nf6zhv
kah0rx2nFWo/Il5xHLeN1lxpOk3ClDcxhWpNGNJSfuoxZAyaraQB5Nf1lp+k/FWsp7gmAu0gJ+td
707OS1i6TTVYz+KId4ZXx3Nmgt39QN3ffhz2Kik9vpmnTyAdarydI1+5ErdgJFRhR2ZbDpaQ+LvY
CZtyubH7Q8HbZPI5f+FlSQs60fMeGAg/5vTPOBU0S1iP/Hj4gQ2s/F6gxnO52EcJl7mQ5SkG+uxI
qqxavW2O+z99zGuIrkJX3d3F8Bvl4y2/YuIiX7xYy6+Mwk/AdWgYXZqYZ3vAX125roK/K1lebuf+
XRUMFWdwJf/V9taXQfgPdgXTwYQm5/eSj93ahiUkWO6zI7nOe8BQMzMLO9tqa2EfVsoISYGKQpNF
NzjYdVyMqCWl9bzls80mDnyYtYPjA0GI2r9QnTsG1iTW1LXvCN/1ce6ka++9jnwWDWeY67LZGTyk
Q3ogUEKIwdT2ONi3sacuUoYNRLNJcpgAqvJx+S3Y9U6xpYLuyfs4dRRZOQsaGAbjBXYV6sPmzJhh
Own+Gy9Bs2YO74LbZ8XoQjfXxkKeLyaLfPOxrvF39pEXAQntV5oGBMJq5rq69vOovQ/j5dmc/o1r
/py0rQ6N9lg51/V5W0GLWaN/G4eM/N9YYG7lKzvDbJG5he3mClRTXJdj8edBLdI0VRKAjhkp5H11
Gb6AmFz+1uincRDy9k+IxsxTDXkTY+HCbplOR8wzRWMQY6hDQqKzak6HBd1cYjOpCKJ8MtPqwQlR
1Dc7wfvzlxR/Gwv4RAgj1Xmbcx6ujG1XNZb3V/XwVHe6vXSMM/9n5X4wyVifgSZ6vMmbyhfxF+s2
Ei6vat9chf6qm82KYUA9BR/lYZpVsPFc4OPPXFBe0SyZOD+Nu8SQezhZgYtrVhNjeoB7iWpj0KC4
d7sS62AL3/a0XGgnf1oQdFOBqH5xD/ncZpnotvd9Vd4+maG6USFLdfDLxw5K+Hko/W/J7mkfsxZk
zntcwiFEvDOKT/PqH6qz+rPping/QUB+z/6mjLmsIalvEiO/7LXRr53URST2Y7kV1ReMi7a6jqc7
jL9jesyKbzTNiTs4depj34E4sJmrIfIz3fg0r7LWJ4EVtvJOtCUbDffmjB6EH/j1AiOdQTI+iVSK
1antj2nCTdVerFqVvS+06AcmWEjz/Ig+3DwTXuh8PmnEIePToJ8FQr64NmeOfbZPKa+mGLUAVcnb
qpaM8HFM2hRqBcTkmzquOZQ8QJJO3/229sckTv79EkjboXsOnQlUMO/nbE0CvWG0sAxhDT8Ss4Zj
+0BuFnaKr00ONlmhxPGJlgjYQHxePpZBVA7LcCapdluBMIYDfBtDb2L1Ospk0wBmdhruu6wrcuUk
ANwAE5fv9IazY9UHWJZg/q5lgMNGTNLxdlCooWjJ0YBTPChpO4gv5RaHD+EqL15p3HN7Mt8/VOIL
sawOv100ZQ7/yuJRX3opKSdFnbDdgkxObmXgc85fM+GjUQIUHwG1H46b7u/VUwOPnehbMUwo0I5e
AuLepoIlFYTqbVHMdIAd4LsAkRrEGg/4osd9uyj3i5kNV8JdY6D35TOICIKP0SOsRsYDh0nGG+JW
bOAwP/HOIX8eRGZ7xUE3qfGgwksfnUtjlp7+XTTXz5NEbm1g7o11klzXqZ3w7nKoVPZGNKjwJKy/
sWlNWjEgrLlPjDqy15J/UYhOUEmU8MMqp53gYkbMnHncdguj8nNbcFJi4zs2ylIhzhdyCQQDgO/7
MNLsUypEFh1v+OZ2V7IKlYsKzqb8acd26qP7eur7q/2a7ulSY/ud2zCXSGRIva1p7S08+ykY22/q
bPSn8fggsR8tY9OL19CyiWwekvTjxoNLH41P3SOWEfTMvBv0FwoQvIDsId+Z70rWQu4m0smmDh6D
ZClfkynWcHxOtU1dtXX8q2gTalk685RrxYtSg7wuB9eS46Hs5kvywPlehJQQD+5QRuPOuITJwhv7
IXbJ4EeRFDMDOEcSF0mZJC/Kvcn8+e7LL91/kTT0piS1qc1mXbz0DNLFFSSwbDLoeDzjS8JDuJe2
/5st7nRqcWMxaN6lXiLmI13+cY+aMC0lnJAt8qLq0XUZ8kDwYKGaF0DiZ1y1XAEc1BK1sZHpdZKK
hNPUiYS0QJ//Dsn5HbsElv7Cfna4b7JcVd95yXbHq07brXVkPUS83wQPCI5V9IID2DEmqAC3jqrx
8p5xTK8QpYSRk538cnHJimuWLLEYmlQauZrQyG4piBoRmGPgWK4+gzmvntku6ZWGLgRJ2mabmksf
+zD1VbcbrDKHJZWdvf5GuesLnKSFVGPdqvEZM4xv8RZX+izHEXR/LYvXOGlH2f5xTChDu56FgeVL
+A+pCV6FLCbK4pIFNdZ2IIhnu9q77m76UT4QlIANBxb7zlWQ9iswryzhilpHQuHVGRgGyiohf1Iv
ACCn6K4MiShV9R9CQK/RMO9/wxhhvu46P4aKg0eAMrSxOgAdbWNBtJLENiYOHv00+KDcaNhsKnDy
OisOuKwTJFihojjelvhSGOrIvmLGroppxY4CDdjsKpZySKvWOu3cDyHRoJNtKPPM6BUnYYzHKBpQ
n2HiE7+GvnRF1FzWwO8vwYZ/zWQLIg+nAtZPt1Yv0nt9HQ83XZjq05CuPi60ChKPP5L3ivA22PvC
GfLQkLJZumUQ2/29e7I/kfVgbNPrZfGDlC+8JcZJW10qhM90FdR7mJuyf7XizEbpdFHraLAti8jA
5Fl2kEZSvwd1heDFOgOlJonAM6NqReYru72/yx0SWcMI5LizH9dTdQVu5ElFoKZCIcTgYOUfHTaP
nDj+JT2zBfuOlv+LegjG+e+x7aylFamPQEig+zCCvmxMwyFRMBYjg7lHkdomTIF6vM/iRAJzHouQ
kqWUASq1dNY7J6n17/S+ORg+gRiMABrQZ4ssb4iHRDTyFrfAM8f+LjGH8uDiLbwIXi6KG4X/ZAvP
qxNvm4T20ze5quYrYu7PAIz6STBkHvZQUZnoGDj3ZNo3AscrPVfOXp5fzdGx0s4k9It3pepIHo8U
lCp6IWqm34Wdy6/5e2CkLB3lXhRG9LTjoN7jgSkWtFspkQWUmrWmRYV9viX1X4cmeE75h2yHvaG4
sW1zfcI591GBS59c25qDtPoqHzgsRzTeSKhD4Y9k/0G6R0VdwRzgeKXWUIaoakbSjQ7w1vlZaetk
VnBBYjVh3dGYqKEAX820oOn35WGmocS20V79pLFLCTOzFKRbHgCGowhgfaJtz/edgXcuyeEBlkno
M3qdGNLZtExDf2s0Mp7TEvEh06jRKkAUFNRQ0CR7OOwQYxis0PW3j6HsUV4wkhTwHZnojzzAlmAN
2fzSW0VVzscjt+CNJT/90Yst8dw4HZ+ECa6xX2Bediz+aqrjr2NyzNoPnP7Zx55A93DFRNivDkxJ
U/q6yrkqBiHcpASytyUqnODpLgiRvhQX19Hv6YvRPk0T3fdCXGshXSZt70VGMq41dUNjPljI/2aX
BTWa4K19ejLAcGjWhpZMnC9+7O+zMVwsyWVGx+csY+rN7uw64BUtFpy1PrsvL0QZtZbiQLizTdWO
kggpHB3Hxf1TrMM4n12f/ocLUMUBHCjsCO0y8ngDupXHHs7KdpxzdxzxhMkkLgs2+/seaFvqe6I2
TzwhNuGiIBhemFnNdWpfaZBYVPIs7wg8FiSeiMFxf/f4lYwimRkSXBY+e0lTQmuDEFLK/jfqQe3h
on6DnyPNBau99KEBKH2HuocHP45/bWxyLDdMEBKwjXovTBXWvoP3xvJvz7qpNf4uyeGIlzETLKgQ
xqFJ88Wzedf0/vJdp+/Drnr0U3z+f2sXyTMLhwtIhF6bnWyKEHKxtThpTWNA/S0/myP6R89DchZN
yYaOG2AUp5nWX/ZVc8qq9kzz0w0qS26PIooIWEoT/Sr0QGDeFKC7EHCzwa17ePqQhBq57jjja2y3
fxwCUOH01dFR9YbMAeoxeuqozNTC7lFI2LCWNHzB+Ryb+ox0WK/4XsKBZ0dLTe51zA7p5rSIsYNB
+X2rMKGiCGketh/G3utUt5lKRZ1+dXUO7O7gVYcYQ/DnYdVYKG4Pl4do94pLVsC25e3Oyrf5nL02
NjNcXrcUWPh7/TrqS10q7H4r1X2PY5GirfbdD8fKc5Uc4gEvk+WP7WH1vAgrETU+uPxhdvIHSr0f
X9ZOEpvqrjffthpmvf7gAZvrnt7TA3zqCE9LonjAYZR9cd+zUSTsJzEu90WVnHu/1pDFlAkrxaXt
kulHYt1EcGo0h6snOlW4muvL08C9EHlnrMbsPkM1NBAKtmxzIHvH48hKH/yeedL1cidHbAPGiA2o
jfEJFYpbshqo1FsLJcD4UnWOBtduIbxOkmP+q9LccMYRU3CwdTTQrYkJ758A1fe1ZyZtQlxF56pC
KaMM2C5beAOFYAwb2Rnq++m9GSf8xm14ji0sJqdnhWHLa4rppLpnUUENRK2j3MQvS5qnIZsUMF3x
ZLzTIgh2IcKS2wB/xwDhG2Js7twVsfgLYz0UtU0aGyeNQn9OzSoNNiKX9Oy5pZxSb0nRo8v92T/1
rS54LegUQtTTSEC4f+MQ7SWzoPep3fIO3hlvdpCNWkwj5oDEDjMIR9NKb/58OyV/hBY4BdEV34PQ
Twd4p/qU9xjHDIaL36C3d93duxoyxziLr20eLixGj3e+EMVV/DgMua7U/02c5Rw24WjIRESqwKk8
e3kFZuzA/zJjLbua8K/kufNnFu4fa7DZvnZwy6zYV/hrqdctT1zPowuCfauFC+u68YXFEn2XwGd1
BnlXk8T80bd50Vxne9ZNXpvmZi9f1S61MW1Tlh+xFyZCxe2ZoBfDF6KXhjx62U1Oj+U8gXrPmjpJ
F+1ouoleR89+3BbJUIwrgeemjr37y57Be3aMTovninSxtGrrN+DMwZaQO11PFM5n+qWnZRikshHW
UnG0hvpqdi7T+IHrkdaITotBbYRxO2zBd7WFjT2XB8s00pl1rX4kZn3a/IDFjj7Oj0Hi7wTaYBAu
4AqWTVXj/vfcA3O6dcKuZLntwvYvbt2sIRYOX7IzpbUYPrTL86GHpIb0lFobNx+MoDP8FBJPC0pO
nYDzLfpDMGTfxr91+zA9eNXHXOxxR/WQ8jGp/wO1GoseHFr/ZUSpqJWqy4TURga5BbJsRMedJUCB
fONVfLzrdQ8Dhwb4sJtmMrNyIsAdhUSxTUgjP7IE/yjnpxgmhvbh2Fpe7572AQzbXLkO91GTiymo
Gh8KeVDvahXXV60CXcqFIaj48jgAyRtIiSFCommBPsDOTAZ/S47h6JBR+RvoMuOvhTz0kQTeTPmS
UHDPntffuW8rdnosjk7Hx5Ohf8q8pM3xCmq2+/6AUdyPV1xaoyOOyXJEC+tULhkM6PPMeQI0RoCQ
OUKjcnVtpb42OfB0WFMEnPosrtfU+/4lZahLMP1mtSlXW3Anw4SVGprrDPtsqI3EdDcHz9dSFtn9
1j2KOsNPORry/xGE5qIi5k+QFXDw2pEm0pI+eNtD9xkg5mbdSaJiiD4liN2cztoy+1Ku8H98HAR5
N9VExhlyjux2vj1dxb9bHw8sD1WS2DFQsdTwgte9uu1/Gf1dirFz+d9+QuqxDTJwOmaaXrqaR2kk
8MUhw3hdqfZIXEjR9vkDGv+j8wghxGCWgfPf5JzmLNz687exoMTjjF1fe9Lup32hgY6M6OrWWXHb
md64tT30MmvFJ5y3lHVc7CpDlw8aCpLcwLTYdyKl+Tfa3WvW7YSyxM7RNMRP7Il6kGL9noaO3Bed
O6YPDpuVii0vgiYjERb7lbh3QachjGe0CxL3872Aq7H73lzQrl0FiiNA/KgVIdNU66afl6bqiB8L
VwtUJrIuaz8ZP6EmO4Ornuj8WDi1X8APW1pOEDzj8GDnPCEpGbGF6HIvOt4X8LZHJTYSK8onH2mH
K1NaQACYs6XIrFq0hSL3bLdM9DbJGELY1sAVZWfQ712aS5Lt96C6NyujCNqv+KHhlo045atXXTNl
aSueh4oe6eiFzXdazSHMReny6D2nr3gf1ISnOrViQ5aJMsbNVOJfuG1M1GCtXYnltdRzNoPBoNdN
g2YAOoouS7ZpQ1LjJFRPiga20+sL+l+Syahutz4tUf03NVuxiJuT4piedKVGUQr0uiQadScYlxBe
tmfRlT7b9Bu82LAmwqA9dfnpxfikwVWc27k9MXsruha/tmp/Q4aCzJF7ifbOc9xlIH+LDxXv2OJJ
ot2FJyhhjuOfZhQ+UvmARgEgVMaZCXDezK91rKArzXU/QXmpqFvQMHNe6+YMvBd7fgB83tqpt6Yh
ROtHuuaoFFX8No7xC+IFDN4UoQbpoX3+u6nt6Aonu/EAcCm2+QBm63oQFbaIhEVwuM5a5PKsEPI7
o5KRx1aVLouvR3DOGpVcpd4L8J/ix4vTWZhYFynsCL4RfsuRUsRihIyz/To6i1Sxvz7YQgXTeGIP
mWYU3edNwTMBpPa9CYBrO9BQpDDIkzczpULVoku0hW6hT7UoMmpENBox8jpat1Z6zMvBGzTG9mpT
Lh5W80nbFpEg5nU0tKG/mi8DO0CgQQwErS7e68iiwirk41ZXm3jljZ6q1R6dnea7Yf1fx1XaTJ3B
1eDF9mXSLq6GMszH8nLWFyXJ1/mcHvDez7TuNBxwH24m02TNphgufm7AucE+u9bgMvbYloFf9dcK
AlO8aM4Hysbg0c/zfQfXKyDEoUqC9Z1mSPowb4R3aJ4w0hg1m3CsNWTpuHQ23IogBHm1+stjC+zj
DJ5thOYK914dF+apDKq7XJWmSvgTxXAv0XvliAjmv3+NRn36ZCibOcivE6Q196Hi7FD8kjwhAOhn
ZmfCz9eJNQbew2nQdCdPZzKL01JjctkAxk4K3EBisduHhrIYDpZ+u/yIcM6+bjX5HovzF39q9v2P
m158IqPZJuJmSml55xyYh0QAEx5QRPJJRoLFLYCX9ljGNmISyRLSVtSSZR7XSInWGSdKPnnA3FxR
5n1pFwiXmW8TqhWg76xx6LdvPcTe2bu5nDo0fKIMzPIeEOm1VkkX6JiO8ww7cTTSHKexvxPtY1fQ
s6bBN/4cnX5fzzfeJ3NxsMyWAqJYhU7ExG1J/Gs4To++/C6z9ffSsLgvPl7pprLuluNfLj5XBmON
WBjWQWGxgVJNiBbdIDo2gSV5mJdMIwA6HwH9yL1v+ZztdAlIo6+8HHXDXzGhhvO6BPz/vI6DD8kM
b/i6FdJZSd60VmG52RtfWeG/6cbOxigZYF1OsMOVHSnpvIOIAhz9eSeSyCHQNAmAGlen475cTeRs
zob+vl3QhCUV9MJidQH0zbKguhNGw+a3xwm6XYTSQhn+McPfLcdfSZlPKoFl0Qo+UUi1apKVwIrd
mOR76fyyrNgoPyzpfKXTKuUco4ifbDkOFzteUOYei+CdLEMcmVtFSw7aZtAoIgDErM3jlY4OLAOL
0gYjTOf8OJ90qke3opQnEJ8Bu5tpCwKNJJMSsp08X9FdDX4XY38RZra4jmmgVzyGxQhLgRrlQv9T
TW/wZOsgA+PLg6svb0m6xVxcC/Iafg5rm5EKQkEjxo5t1ivvf2tD/jtKlTLL6HP+2/gE8PWB3wBR
XeHye5q3o1FH6JFB2kqnVaA4WeLszze1JXa0bp4sFjscdOIoJm0RPyZ/+tm4o7QKU9vyvPJ8Hagp
E61DQjUiWl4YUcvBuEsdyKUGnkoNDAGiEwzuXqeTaDBEXKRVF6JpQIUPU6LzMAixX8EIzLCXnp4l
rW/fZnp+9HrOqqrQQevLiLw5ZBUYW0OCLxbJQgLKgjnP316BffW9KIQLcoRfrQwLiRR1/+yClC6e
4hcH3OU4HFXx7yfSxAsw8sS1A/QiOgb6sHV1GUwH95ro+ynxguBnk5qrvDy/V4BzJhwag79PnAMa
kHumJJseGBlFyq76a4iucvB9VoyYCEuhkNrMBlQkS+lLr9gKuO78K6ggWUXQdDxmyIxtHoThtAkS
QmAmmCQjwBLIWGtWwvp1X2meTxj2Dpo6HA0XP1cJFnPcup1ckS199k8TnOvuT9lKrkcA5dO3HAjV
isShz0gfyImexGLWKJxjx8nic9gq69A3MbkVBDGYH9rSSH/bi33M1HKOmj3pwUre7Ruv2VbZolD1
3iopg18sTg8YG3Odr41CtLblh4XQhvI3XKzbiQZ1EI6vOprm6oIDpArXVr+nNqYSlOYU358/1nOj
WVyJgbqN17FUayjkzS9/HebkT/gx0rDEWxZhngDd0wbrKv+SWt2fvldl6J6/mI65hsVjVqdOr/iK
o9wvQS5q14GKt6KGV7jERvgHNajr3QZpVbAga7uzK3yQkb63Icz8hAp3PPZTKMr+688PnYw5gV/Q
xVLXTY9HlqHl+zHZvMl1dm0KrRYril4HHOUpjFLUgxPPu2yrAdkO46eMl/rrq6KqrCMakCwP/p6Q
dViEO5V4o9sXXy59rKA0JszsJQOFAe/HI9O/8xC/xOAqlvgXLLGs0t+E4oi3DoAHa0cT1bfTRUF7
9wCwPMIWoqYH+7q2KQbJTZDH37PBBCPBccUnw+7qilSiSFM5/kUYkiyas8AgOHJ6vYWqeLSQNyvd
/wQyWe8ty44ssIQgrrSQmtIGA/wD0d2Y/bsM6B18W3Hj/dO9+jnlEc7m6tqfLFWfPpINc7PJ23Mj
Nj9olLUsn5XIuDPUuoLlKuEjQpVQlelxNSluCJuxCdanK2hqd35l3yB6M6Jl/P6qLxp7nt30HD5j
D3+owGs6CfL/sQ+Cw4zU1AU6Q9q7QGJCWOVqD/djTEs/gMdj4WbkZTVk8iJbEzBfmWYVoKa+4Y3L
vqmmCH9graIj5fIi/1D2Gktl1J+s5OJWTIhuCHWBJPJEUNHDxZfvF+kYDB0i8bGyV8jJOhzfYpfy
lkx0TQ6g5Lh5PsPaXFC0sFYLBl72IlzuiYKgaiEldEpINAXiYbFePiovCvoKJ17EyBGxgl+FbRHf
eadjnavXiCHKxYGoAdQegSv31DOSxerGNzYGtz+ryCiUDNjdwKiU3IHqxzvCbQr1h1CAHOcfvvaq
aSPs3Dpz3yGNMr1HNJCIAIOIXpRkEYrK6Ncfh0mtbqnJ+SwDNIOGrt7GRTw85NWBa1h/FLeLY4mR
yvz7qzdTwjQnIagZ5PKoD6D7QEavb8WyVK82lzp/X3sTlsh6UNvc77XpWY6NJXTCj4yXmNqUuI3e
ojZzd2z34pjDyTVSdqziWYOiEXJtN4jxj3QhWP2kQMxwcSQEoiLfKxt19Qe5GfXegdyO9nhczTvO
d8k2DEZvzOZ1xWNYSoECQJ4FLbruOx0f9SrvMYFNUlazbwqa5K048HVBXvmv4NGlfgnBXMSMdrub
eaD6ZvoRdjFF0R8bEREfpMhJRzKJUjWJ8F4PqsPzfbsf1taklH9zm5oMnpcK7Q9LQ5vea2uUfDL7
/GfoYTJzZIXwQLVysHlH4GEZEnKtXnoinqoFWC+dzyslxPuilZgI/Y8vnRUiKqjDPmtJAE7VwpJq
XyK3Y62rbJtzCJciGAbrpWNfgrb4Wyrv/kEEeYaxoMx62cGd2qSXIL5HUsr0bK6GPzFMb26mV7Ia
Jr3gJkgXu2C8XDfSxonS301Ki6oz7VGLlDz1SgxiDVdqGd5fA2T7J2IpQ7yebZJylPvwcH9TyRFD
kVWDVOBseGeSICJotvAMZydLI5bM7DV7KM07Ns+I9HBJP1bcwz7CjW3eZ3uj35y4l5lnOdpaqIiJ
68fmqVm4lr6T5eEhmr7HuKzikaA8DudAAzTPpTNYvugHNZwvFuWZVRBYGyuTOi7kvHJQFQMP42vs
dVt6WOMIBJ5o1ydnT7CCiJFroUUBEKADfElC6+P7Zh6v35RRvqI/H7LYwoLsuH62loNWG9eZTUww
bZ0b5mo1Tz/DdJtQ0PBp11xYMeDy+kAo22/OzN4F9KUlgskt4DiIfJZU/8puMIoghkecKY02ULEO
6lZZ1ZRJUJkM3/Uu3E3VdBPDBeMLnxHR6hJeASfpdfnnYqxCU69X6uNeKmUP51QmMMV2m/cJYgOx
ZVnQ6/hDzRxMN4ckuOtEREkYQLaMkDmlJs4rQW1KOV706HLZtux8kVyyUnd8+20wo696nHVbDvQZ
YVL06uhgWYYk3ZxZUjmUoeGwoU0nWvYnx4VoZb0ClxEJWmesluEIlzWY3FB+S65dPAo692idesnS
ndOkPqjyuvrAN9GfBVv2ARF0SzRGV2igxKd90/ALBHyeqQuyvmC38sUU+Jv9a5w3W3KB53VVBOy2
B6BKCT1PaSNZq/+6tK0j5H/7GlTA3Hoh/x0JOHz1bgQdx/XOzhA7+81HF8WaZ4oyQaxWfskIM4Sd
nelOy/QGdmd9hMkwPFNgMJOuhQeQ0BECPf0GivEZ4vsAUbVt7wnuibN+yv1zPb6qNQIy70/JaRoJ
PQ1ogI+bkDKlumZj/FrTzWSY5KoNu94PteIpAYGFpoXRMy3U0ItOqbtlFlkz4RRgxtceSbK908zk
qt7+hwSwVav39kuc98VJD7oH3MyG64lhHIM8jE6kaBVLA+y+pKrvjGwoV/4mS1EgVZJcxyEpTnOE
bCAce0NxG8DxNqESlxumz+A0hxsmQKnMUj0DbgwItO/pFOIIhmILBnvkNhORtxaQ2RATJcIwMAqf
5vBpaP/uOp2nV5mplwWK0J4I15TiHjCxkTCR2lme7Q7eZXIeqgqqZc3QYEpZXjx18+Zb3L0MoBjA
+n0tiFb7FF7Ot/bP84vB6KoLlv4Ts0zcO23UFg5kzB7ZUvqc/pcIAaBAtqgcWjQWqy0GJ7jrajX4
7dlBLCcOhpazwZj+g0tYxBGmfUwvsXYxOMOHOnUtbUQPXtWlw3d6txQynYvDWskqVAmwZLiZ//z/
XKn8Xa5MWXMsfOs0PsfsF5xatowB34DB7oyqaMW7CLfLFcjHy2EVPZG5FI9y27wcVccHgtPgEvNC
4ug/7+ZcaFmII8/Ivs2n/aRqKkPPlIIpoz4n5JZlsUMG0TQaCctCFjM42gdrPDjU59Ql3o6Rq+wC
K4hJcvTcBjwLJxZ3lF7qLYnyUbNcKbtTh4YfumzSUsn7K5t7GlE7/vFC0hfjr3uS5PLv60O4woso
xUZ7zF4eFay3oV1QlVwSqs+mGZASXmtHPpwpIJ0knlpv8w6D9T0ENKWV+OKpJuuCTW81gSbbI0XI
bMyr0/LMvrIT8SYpu+Q+9jqrB+VVUzcskB0202eKusymW4RlLjvlYwUUsFMG2SY5fzRP8pn+GfsZ
hEa6KOIzFApP3+zVrJxzK3jtwWrq+IyM7UbaPD5BKlab3RIfGlzJ26c3vaF06aKWkZQtRbxAJfQI
GRjSY38vADJYnkI73ff5Ifw+3/SZgsF0s4wOkv1l8cMHse/9PAi3a39cQqqXWZel6hs/kSVU1Tfi
xW1sJtpa0ovP6OK7w84HbI0wQV2ydYOnPrRCP7puoN5jOt1ExtledFOZkWeyPzc67a1Bnh/jNNHE
zk4atP5IVJX9SYQXENWsCSXhIh0XliIygZH081zTAYr3oB1VtufVvlOy9o4AeFrI+dfr26oRTJ9m
k9TGIrSXQNm+zMxZP+Ja+AMRv0s9nU88nCvLd3F3HAuvpYtA7ZXJGl5Y3bmKkgtsOUWpPSP5qlO0
LHJls/78C2VaKtBEGvsD0QjmGzPJyiEPI4ayu8xfT7rxdKWMP9I2w6Dsy7F1k8JirW33F8wWA9cT
W3ZBDF3MPFC3UElnxHMtKJ4a98CbXqTsjnlivGaeqs4Qqqih68eP5UIc7fJrDD2eYF8+Qf/zTUDo
/ZzZUdkW5eXtYczcv72+xx+oZTKw+EZrrxf2DtIXxVbwKkcR1vaQDdxbAxudYNdLl5i/EaqOUfxQ
i+7HmtexAxSAHAv6jYRx/Xx62ED4v4KX4xa2Ln2gxwhyFebX290Pock21W4b9lZKnMTQgKekGeH1
CpnI1PaIgGBGZ8HGM2Inj0T/boAJx/XwU8+V+RIzKn4S/2n1nsf2Cqzyz8icxoPrSgfWd9Lyht/8
LvM0dNJlPrvdnEw/c6tIhoPK1+sxg9S4od4ipSHVTukfg5/bDtnXggYtL2Ie5Og7k5WW15an1Ylr
8AH0sGivlVdZrO7mqjRUSstEhEiT5x7cGA8HOyIwOzlqns/Pk4vNonfbKmoIP85FOehTe5JkwlLl
yUYxA1LmXr5yYy0zyvd53tmB+Qs0mGZQdm51FWnfoMlsaDig+gLyJo7PgPGT2IvMdTBWgpYB5FpA
o6DraTbCV/ZjvDda6PG/7d7eo6PRJPgnkzoBQUJfdsbJ64mMgD/VU4MLthn6SYUIwSzBedRKHyWJ
gHmjp6JdMQoXzEmlF+Z+yWhDLkZTir2Zod882rrHkIecL++2ewWQVuIq18L881PCEVkCywCuVFi5
hYAuByjiJRczyW7HFceX5H2m4UFiqE15F2cw8jLRNWEFb5PRscnyHv0C0OoR45nsyh0ZpQ9Uaop0
v5Tnhm9VbUhYGBh9QK+28ZsYvmlzH81EOLnEQB58ReQZ9VNl/pLDkFIPcEpPaW5aauR8x5mlssfT
g1Z+TSatiYA7AUUnDK+7FpEsGbh9L+INgPg2uAnt4vl3xC56ZFuvRvdJX/gGxzYw5MWOdPVRrc2c
aVLwhkTbFMygsBrHktK8BrxTwuN6ZAlJ6HflvpVZwArhpz2pH3AxO4FWYg7ViYMM0bpWWdRn2nEA
Sl37TdF8NK4t4IlJTOw6SygDr5Db87h5WPR5MyUGO38DIZA2hy13SeiW1dOJq/AAQCNTe5VmsPqK
B6YZmnuHIheW9t4MDs7hqXJgmbif57PGxgXyVLN2wYkCwsT8G39sSUPpxcIRTD/sf99YmOBheJeT
ulc+8C6frtCby6ZyrRTlhAxv3Buc24ueEtYAG/aZ1z3uEQ91ovvi56CrzR8uXf8+SQ5oI0feKSe2
qwOgJ9QCOWbp3CeQ/gCGVOIHkJPCR7HTKUqfJalCGoLv03xh3XpLK3/tId7eqgWNY7WCvFii/3Qh
FclF2Dtg12v1KbOKQzt2KZMDhrRNVFLupq7V9oJtPGvra0ndEZi/KjEBvAvglNLmVjww52qNKjel
2D+zBYrydspLksR/4yIoPYsd7T5r3cPag5g0qrD3NTJUJ2KS4xOKAgp9TKXJWk5Ogj3un47BHpvt
oVi0M62lNa/g34c9l0Ewp1uPcpD+4o7Tn3hisHUk0+LEDhnWqIqR+Aim5WCRmXzzAdh1XPIE6/9u
s+1Y0abt5oQ3VJb6BIpy5DED+XtQQZaR17qa74VIvB2p7nJRD+uL+0cF4DZGIgmnXrJpDkkdPvta
1JbQ38X7Fe2o8qiDEZ7owAdDVqzgrfwN73jc7l3TDgC6ATRrC8vJRf5AiFAKZvlPmx1uiQ6dAa+5
5DPSrESUBHbtOCzzsnAfnLYoV+olTUYv/2Ylbc3fANHioflYwLfx/57Th4sJI0QAQoPk5sZYJNYo
iJa6gHD9BkqfPU9S8Vl3nAYLQrScvgTVxgm+Uhiq0Rk+8JBut/YHL9i0wxm5Xn0zUJZ5XG7CNei+
r25wK+6u9wt4H+EbdGBbdmcjUkp/fTsm3Lobkz1yr7x0oso/PAy+u4f+UJ0JzuSrerdKzcbJlOdL
+TWkuBgmINdK4b6LOw4LkWm9t2bxQtXahgZaMmUBeFqG7mwccDE9MkDTZ7jOYDb3cfFtzaqmvF3j
2y5aAYDFwk3wj1zDZqttIFq2jsRcKJIsN1gEpkKA6RKieJbOjzCFRXvaIgMjxMk8GEHI3JTzGpXu
6/r+KVyeKVvFWmIOMv29J4ar5aux12W7lVl2miy+N5UOzUNublRO5GysCtt7aJi9wgfX4xbMaGD8
MFGNUj/ie3BbydzFW/MtQsTs1R0SwjkrLw34xCC62C2KBasy+leLtXaIjtC6RuApKkpQfB/EHxYq
wT7AenDg4xH5uOV9T5i2OsSlJOH/INtb6PUen6TQab/B2/MALNERykjHMMUr97FjjdQDTqbAe8SR
//eOJm4lRepTrGqW+kCtemscdJYEkdPKwYLTxjwl18d3aqX58ulbE3gfCyLJS+BOlriw/DIDetDp
tnmsZKljJ7h8HY+jOj077AgePmA0ACEDgSzd4ty2EfChX/asGxJIBmfysWtiwXCDdymf1v1KQPjt
xVZZv0x2rhcC0dr8jLHO6crQCoWQIXK1QrbfU0Zk5XpD5koR4zM8b78H3vqShhCGiqX2LuGFj+S0
YIH9AnCbXYMGDYpl5359HSz3O3bvIlCus+sKifF43kij3E2zTyypGaD6WLFYCIFy/I2sJHCw9j/X
M/kwOJFg2Ocy9TV3TBzx79LayQ1nuVCYhZ/aTT981gCXfcbDKgP+ocZejeocwVE1yCTO6sDvD618
w/ufTzzDLK5Mc43O4VCaf0kWuN6u3eMOGgeI4la7eF5YRNeqoc4kPGwa35QBr+PJ9FNFRyoW+Jcn
f6+q3Aem9TrOrsB+jO88oQZ2vMl6vRPj+h9+6aLgF9EU/oEBECrS6PQyuhzBreTsi++ppkKkpwAS
WukIx5dc0H4sBGb0fKBJd+G02QJ0m/BqUrGiYr/sga1wL/30OQd5Q+q0/FzSKrZx6TimILnU5tnN
Bu33uHckkfcdankvj7D995hei6tTPN6lt2dnpYpm0a8RzGHiy9yluPScURmMxxPYvc1l4P/+Uz9b
18wJGrNDb/lkAFPyu2/TkNu6LY9uT4crCy2dax9/CPgadzfwT/9oQ2vTgylRIndBVGXkL0hXHtfb
1YSgXTIX63fala+CCzo+dSVBsm7S8wyoUnVK47UflRIrpHFXJVaEw9C0iAghpD7e8+KpE9hiL9ra
jruVXbppEthYkhoHTN1CrCsnPELzAsbakxC+T9FrFjw7UFD9LylgDDgfsL4dDISpOkcmiUwTydQT
0O9tzowBO4dFBIfeBRV6VZVrX9/i7YghB9Xe7M14IbjNvFtnI/S243enTXn3PvngSTnUTl0YX1+E
buMk5j91qEcOAsqpKi+RDV4FjgnF7K5XD9tJ3xsV7mVgjF7Vnv8jUJyf9KmwVR7WDEbYE3Wpc5FO
HP2BPtMX84PbNc0GD5sc8j1k98uGNIpVqzLDs/F7QCmfBXc8AqRYwl2vL1wVETEwztvdLgeMf1zF
OKkoa6pMo1HoVwf1FWe+r0SKAAR6bQSN5hi9mQ6XSjsHWzdkT/Py7BiwIR8M5rUWNzgVRxFepBKp
W2Q3C+FNpUuiOqgaQVNmdGsDQSpNPVwDa1JDYt5zt37CgQCRYgRRrsdH1IqAhsqmGCKsbqOIJHQL
8qu6/Iqr+Z9ULTO143MyvZsM5mj+3KlbivYSJfK2C2LctGNIJFLIW+bNqt22BIrXL0oVmxoWNkDY
+/wurjFbtIGER367jZoZeaVL909t0wfGPrgw+914riO9eHrr8p7a/Grf8UqiotADvl6A0Tn5oyU1
aNWi+DN/uBM0sNI+Gu6JiXjvs1COUlhmdgRcAtfEhRGGCTYBbA+gnVXxXvrNa+qIM9umK1005pVF
b6w/2Gi3XmsZuCb33E/5IRVzV9r0djfgIDUcuAnkZ803Rdhb9mMo6TC+DEfeqBZfu+N2YJZNOZi7
G/KybjWZN0f1zxigbc/4Dfi8SZrcOaFLfpFsvcvlvD7IBgTCpTCnxGhbgsBWLwjqrF6dQivIn4zt
9WzmHk1n96MtoPQ64usErq3lYu/+d8GF5NsHkVh+0HYa+nhWWLS1A8dvC4bX1DtbN8fpHOeE/nNi
lon6UYZ8tuU0dRrI/9iNHwJ6+8BjlljIFzbiuj0BcAmqVKsq2k7J/0e62MR8cj1wyND49Hr4SWh4
sHNIj+nSkD8HzEgZbZ3JNf0JV+BgDNi/7AEhytQy8s+aT6SkLc8/XsfBcU7+Wb9W8NdYfEXouXsZ
9M7pxGCKnP8k+asOO1Lb/rXkAy4yYuCpZ3woCMufjuHTR/lwJJxSPUtInbyKLM6Mcq9pDqFIAzEE
6pmOwvaMf3Ynlggh2DOShiOjIPJsS98lyytWuH+T+5bPVjtEwJ7h8QSkwDhG8pxnZN946Z+b49Kn
HHy/Kub7cSIXszM7dgplTpiA9Nc2kLbcVUIoxBJfW4SIOnjQGfAUiyVVV/IhBoXKsk5VsBV6d1E9
dKxJ94UXZXbcNjjTfSPjckQbxs9wo6nmtKH5JtOT3Iif9oI+w365Q3NLezY5YYZhscM6Ru7WDOnn
dIGxE92mQCWtC+LOi2JljfffBfLdkV87AVm3MmGz0+1r8qlJyODhZp/otDCMo9vQSBhMmNbQvR9m
i5nZUaDH4H9Tvsjx1VJ+kUUzcSqSoPvYWx6zn7Q2obRf2wgBOqgSc+l6pmwZVADGEELy17HyEKvv
EODgNxJBZWwnSs2EUL5qC7fb2x/xDYtmOkq92oZ8OSR74i9ffO1cY9Ec5IuLE2wEwmhlLjdec37T
ZcLkdDJmvgpmrPKW2ZH7AbG3DbEM4NeLuOknUyoz4OckBlTxGpvuUWsc9iDz3wx7dqKEcvm5g2N4
EWU+cjAJLn4fv7sJ3rTGeeW6Lf4QsykIcy4bcG7HYWgdjKRW6Ij7S4KPXUG5j7UqLkkZIi/ZInJA
FhXYFNt6fhZljnB1RcuqTSmFa/P58+2vFFtzlNFzpKD6E+VRyyTfgJc0FL9WN2jYUtbOV5sSBgT0
zkisvIHwMtHrDiSzhOpUwKPQhZ4XM8zOVLD/Sglf3f1AIiqh4zS9ByxMZjZpFgc8dAse0PgLkS5K
vg9ySSCuJvA6Vbt67t2nzk6Ab4Uc/WxcQD/yofsGqyzi7JxdHSSmDACwuyFDLThWiSRbEvXNXEsk
IrX0SwCW2XomPDjvuTQf/w9Hn0HdqqYX9+SvEbYEVqOev7uKSdRWbmwttSaeziH7rRwoDAq8FGNR
AetEGlINaqt26fW2wBNL9hjG/7KkdjBEAJIbb35Q+yR5GIysZdDemBgZeoYweS9xm2jWPeR/bQ2C
VFQE3Zwvcwm826QqvrvoAaPyX8NU/s+u20YONGqYD1Q0PNieAQu49wP4lAP9TwbShsNQxd53LpE7
banD8Flm9atoaXcESMTbnhzdqhTOVeW29zsd7H+mHERirWWtA969ftioHSS9CriTbkIRXkssvfgx
zXMoCV8vj8X1HNEM4ncP5yNiITz4A7C+XDg2u7aKGQr3PP2fv5ChnQkhaB5ww1CA0ApqIIyPW13K
gWxCaeHNEjBxvx221FJGxcHyb3TrApznGZjNsWNr4AEuOAjod1tu10qf7V/2bzr3QyUAubmzjClk
VNrj2n2lyj/qIKrgIlyo9GRzYnAKIqtOH+SJy1+JFKpeUfIkaDE2JNsvTVfD1pEu2h6ljz97bIxP
RODolm29WbsyqtK+PbmVLSr/43d1siC5jpsOpDZZARFoch+GXbh30HBp3T6HjeqRzh3D0KUUPvRm
Ai5ox7V6Ip/i59z65AXlj/LaWRjBVTIpZ1lqnEVYfaAX4f1zK93EQII39q8Z2Qm91LeyGbeVPx7f
xuEo+QUsJHLlN1cb2n4lcrU5x8W6IYpZHJTufBYkK5rl1GlhuYN+tXUbodrb2G6eV6gxsDjT93wn
2xmHEzMmD3U8wJL358Ktude7OBmYbxsB1gS598rgnhVH+0QDvf/+fqIM9tEk8FLjCTjVQ2ClLIVD
d9PECj5Xdjw7MWa/FIRwCeMwlJNp0aygYI073Biy0cPMZPFgBLiFru9/E4Nn36pBwGT9tFJfzGyK
VTmO4WTL7bMD5YiBhR7fzsWGeRaZS/TjmoerOudNtAzM5d+pRgD5s25JlH9MZ+vPyGR1LgAlCvYo
NpxussSJFqj87Ij2rJFzbCR7Tt4uUqkWY92jDJ1/9qB4xW/0NK2TacdJAs3MpRCKHd/O7EE8MYP8
yyqGFO03E+Thw5bKeYmx83LYpACCVSHKHovogPvm+wlncAYmgdExx0bRZpwDJQauPkZWE/H6mmMP
1Bcw1CbN9aJ2sffzt2YT/1scMryR8fS2v36D0++sS1hc+EW3kdzjP79LEEgh21QpvsgShIY1plBw
uXSHhsCBY+l4JTklw6xJnSrrcsVNfYMlAku68m/97KtYIJiefaWcpmmxMww6fD3gtvxQwQ7+tzRD
dAaI130RHOFqBXROK3ZZa4IS6JJFpNwKSVBFPhT0F6DKv8JjUVLgWXOuJnNmOfiYFvP/xl+2sY3O
pP7iwJrnur9e7UPqt5qehpnDoHB6fWA6+fqurLFFlDreY+TzmPYcNrv4sx8aJUv3dWrz8UrCyxv6
p9007zYukzwxO1tBU9/lZwXtMs5rI86QP6i1fAnHRdNX4GIcR3/ihdlpQ33y/V+TqdpQx9FSgIz8
Q7qKpoVgndpCV8jJi3YugaFJJjy7keD3+WgRVKM5HYoHQzohlwfR/aGTa6FEbfjBPiafXPEYT7wN
K0uwKcA6GVmQYQMZnYEAqyuh4YmGqWzefqCwTSRU4QBYDNraiSrlNSgBKc6bNcaN9HjGVG2yDDdL
xkN367eS/8iNlgDWqwplEk5/kRF7q0p4qfJ2Ggmw/yFWrAxNhHPznRrUb32YsMZG/grdx/ebuaD2
m46h70ILq/EeYyVglIx9UM4pR+betyHE4dDD2RDW/0Ugur6flGrHPAiNN5qAjx/p8vFJiSKaQqka
3WYOpzazgk8DLJToA5LOBGd+cklYa6OEq1WpLCrmpmVnEkGpo6m5Mt5THR8WKrvYGJGgwIyejXMh
46MAfIKXuBgux6Ybk4J6lylF+8jNr2LBULZVBN5dRP0/V4D4D4eKCHXRKJrg9kJ6bLhfk2iuJa6T
xckx7vaJlULCLcAlXNihQ/aFy5XU4ydHxmnmx7BD6+8JEeA+kKI1OKeZE32bQ5frOJSECOcr0HuQ
sS59uIiawX9UMguzSSiRONuvM/c5DwZ6KMdBEnkuarodCDMD8dm+FPBLQJB2Es8uiVYh+nuvwAva
2CZ4W3RO0S5RscuW0xEYA6f0ZDnrJN1RXQ4x1bUD1MYGrA1vnESolaWDTqGKthQNA16u8zVw5I8a
Qa7N5mLstAwHzskyzwM4LrD2W2VaAhZqUdnhvOVuwlRUD6aDLR9GZBE7niPIGB3sOVQ/BoV+Kkep
Y22A4BE0wN62XzrK3Paoi+vDn1V01JXEXb6xuW2MZAsg8mJqQUrgu8HagdEhootRH4S0cPtolrOC
ezOznkXQwxD5OhQ2P/ZijWaUBbBx7ULyGjIqPNs2gUydNyvuXlrUv40h/9POAyIHaH7JI3ivNurR
ek9Ri5AFSxIaA71whQShQZ2XLjbI98Ig2CphhNvENCNLbkTRYvjzQXPuokF4IuKAe++sVuUeFWhZ
xdRJ/EQxF5mTtzI9eHlXP7eSc5TRX/xfCDeLIKbStjsWo8LAOBi63ZZbtN4F2dmouvoniQNRsuTX
0tAwBwQLvmsTJMVPGsOnd42+kug7d2qTQ+s4O7Ltogy821HCC2TYRpNO+dCkkFvq88KWgXlNmyCW
Yhzu86uWuG2EppJiW1F91cgzIuk5sqloy/TllGyptO9wO9O3+nO6ZbjEfwLlCGLO02G5bxdeaMWY
4pynd3a1hNztW+qwhzsX28TtsjPFVCa2c2pbzkCTkQKUhtRiQfKtCoBKoD04Rx3Aj+lM3ZzD4J4y
BbMyTMV8cwp1fmeKmtCdBcq0fFkwSsEYGAMNfHo7TOkcY/AfEiA5S+wO3qCWiCXTqpP3+nHbPm7s
WOmfE5LiLzKpaOwe5sQcsUoMBRyPg0FhulT0l5bqGpIWUynfYtwtcq+VW/BrCAjQVd8fqO7FmK/V
n2Ri0f5H1b7by7JsRlpz8yxRrwtdeddSF6Zf4B9Hxu5ZQXrWiPvu79eCvcyhm9F/v5MqRD4XmEzH
d8RUIU1bqVVaapEAYMg7owIOU3Mxq6nbkWDRjFXNBskxdeK/EVLVf9FECff1270B2X2RYGipzFT0
ve1L5iqodOVczcNvLh9++ByxXf5q5fs8Zu3P/vNO2Zo4U7GB4jdkjM7L28AS7hmhm/OovvUj9K68
JW+Hom1Zx6n4tfOrLnaimLppw1J4BiIZdjgiHoTK4KjVdg6Q5yv3bDLvRlSuSFY74f5bsk9drwdv
OWKxGBL48vDQTdc8azRkbn3v8Z6UHcZi3HILHZ6WgJ+4RXLf/7rcz4aTAEX6ZvGbBwrKqak/PvJY
lHZHedsClG+D2D5uiUKo1gNQsWloxJhRod1W62GWvDIezhIAp5WIUYckZCJ3PPKVgMKdoZZuHAor
p5gqSrQ/9zbwQ3DzT/YSYJBsRyVR9Mc3gN/JFBmVTxb2lwQX64oUUV27Gk+RwltQRn7HQ5gUDoQq
DKE0ZgEWvdR2zoqiOI+z+ifd571lMLy/gnAnUagWCIVuLz3FqOvy9J9NncSwU1iVfSt5GKkNy34G
7tcL1gDdCQhwffJn259yLSYzowk2RS156G0UTlGJSLlkwCc5jbHAoWE/V2YTzzjSP4HhwoJsxnj/
BenHRYPL5baTbFX82ySJAILN66pI2lu69UAH43A1PXfAI7dp4wGlFwkig79AZ8LCi6AcQH0QYYsq
V0sKYrY2agnGzBlAgklLALhknJHFq2QEkjpwkPV1M8NJ1oShZLfh5llyHwadbKfZejQUKd6f11zG
rKQvfBAul85gSJq3tk4n/dc5vDQ0BECKRazwVKgZgDnqZ9yZi8dbgFjaxqIgfItgOzvc8qwRc2ty
PeoguuoGbqSenMXjLjKkDz5MXr2r3DaJSjbbqgPhF4BJDdmKYNwpONmCCqcBioQjuSfk1cKshU1u
nTl4H8lW/NU3+waIEQFPja3EBFP1TBjD8wvSqRMhzp22weTeFAJA3WhAsmAGOSbo0iCZ95kFXnj/
PL07DMtBtV7FtIpLlRfdqFZ7rENJq+ZTEy0bjrbgJzQecUK0ybCFA8GsVS+L9Gzy0Yf0KJeXFZq4
hFfgQ2P5qDlEOuDxGHssqtIrW/2NFvNKA8b4tCB0BbJjeOYW8dWhanQZcvqJzF3s3D/xXAcdDAXl
f1D4H147tQwH9j+a5W2s/oFHdDooUQ44CzI/zc/9p2gGsSIOLpfcRuTy2QquZFbX1v6x7mKADx8/
mQq7u7571dUYpUe7Jh/ufD8bZ+/d5xHL8k7oLkJz+eqfg53mwLFWX2NKneyTn4GPp12rH8M7CV9S
orIfSSnrq9kg2xMLqKsV/zBC/8CrP4/9z/fmtDzC0fJrPlhjrcr0r2j2Nx13wo1ZxtMuuR2CRZ4h
42mtQUpkH76ePN7wYZf21A72LFbY3BKKBmMt08H7i6Du7sC8OuJfqn1JdL2NQNmamF13uZ18ar+l
Dab5OAx9iNLM94QqnWkauKFgJlK3gmW9Me8eAeGNutjCNb87nXmHk6VMZ6tjAyx+i8BZ865faWMO
5rpAmi6/jcDAC988GQAXMwuxaJUVgaVge1hEJqC1d10ds/8LPbcNntib0S8L7EjE8WP8rvbate+L
4EEc+1eF+p8gaU6T63ytr9oW9dmv7IMIdX5emOfwK4PIwTutXAwvy62TZ6FSc9v2m6gtM/Dvh55E
Pe8/uxPl4xbrnCnp5OFL7T4aKPRVrlA8UeLFMvsu3AWdeRusFyGDAudJB7NA66Ftj17FohwWCo88
yPPntE2jMyyJzumscaeBqC6+GHTrmF6u7+K4RNr2uwsTfN8SOhOxNK8nSxxSTC44lFkK38oz8oDW
5gOm401FSp1UHrtcx6Tz2NRfAPHQ0/Di9Yw4sXo8fY03zTpBWPpt3Zow5zWbwCCItE+VUCQBgA5s
JcmeUaYZWJ0LMVhPqhdtlhfNnui3aF/VIE8ANXng4N5TLZReyRaDVvan+3mhDqbH7pNa7zvz0Oy5
kRCKMZQ6OBYJJyCHxtXq+kfqVjt/rOckU0qR7u7537+BfecWmTKY4+fggyJutSDehvNzIpsovlKc
jthaDXmKm53KDQUERgHllaY3ThUVb9eWnTIqI7fNE00SG6jlwE9rvELSiNK4ubNYWM20+NCyJlo+
gfk8P0MhsTqjf9o60S43LuVBb/n28/V9p6QK+87dTyRvlHKHRTCfoRHoTiIAKfsHN6hwZrzVgToM
DMQ8EepersY2reIq++hcgBfcpM8K8mdPXkwLTtwYJuEragyZ7vfJ+XKcfW4HEsaF27rabw78c6S3
FkbL5VRPaATY/A4EPWVDq8SCxiOvk+8bFVW8xpt7zIxmPriVQ6Y6A9MKgupZcugI4V9gx76ewQPA
oHBM149Nd78iu0v7uSacYTjSASnd1yn4e14JFNhklsNY5EZCBe8WRmL1GIGxkF8Zsplk/ev5s+ty
IJQRcaJ+S2NEbZJuOrps7Bo7sAiYjD3LagYuDHKc2VoOxH7o0/WRB+uHgQKEnLoQvYBwvW+9MF1A
plswWaw9WGc1ez4hmgcyLRYnA0Ajg9INEUpf79wrFixzVT0kA0dg52wLVpg7KB5gOG3+dcJ/0EmO
9FvFSJc6jEyAWZVe9TCaiMdLs967+GIw8K1l7OB+b39TVm4K8rcSX7hPp3pDEdYUeHc5OZEKmVwu
KU0m4P2/OLfzYmltJ6g/w2h/r6M4bNWXaEXLNyxQPy9Wm0bzrw5/B7itEmTpDj8+7sT6ZPW1rRl/
kwhm3x9rWfy929PKG2o07HgBrd3JJjBfrxXQbtcuj1wquFpwEMndOQZshfom5LnuM7UUMhdNzLsM
IBDyXwIJ4ri5bII8NergIBWzFRv1/18HrFhcCpkRaooQEyqc1ok2u9x8gLu2mZJWTdmfiYLi3NnO
7ocNuipmfIG4mQwUffTQLLoFsovZ8eMsEb52HCTfT/0pJLwgjKUEiE3CvTRSS7PgrIM2skNsKLpi
9UKdGwy38hPbA6N3kX1eqxRF0s1A094a0ZjaOZ7bm23S/HdgZOdTQBpVaxFEOfLnHzAdiMzp9rI3
NLOAWLO23T1iGRCkqVGjNTG5qjDGZ4VzUWAV3S2sqqWPEjHW3zL0frZt2O8XmDkFViphKEykX+6+
fjzR1TZ9F7+LfvaPig8WN82sGpzsV/lIy94vy+0ApwQrPR1fbVI6D6nOWx6qXsPEVZM77Y7rHx8i
8mTkbC4g8KfqReywOkvgTRTVVxYB3csPDdrPOPHfD3pdmVXEwHGjECe2kQ9nnEQSOaZha4np2GXn
inEkNgEvNkk9PMsZhRaJCYMWy1+rMR8tQZNxs6bNsvUjFtcIDNI5kXienYO0XRGlYPVKDW0a5kPi
RAuE+ojW8oPsUFkPLx50bNZVIPkPAQyaykeO2kcaM38lE6kynmZq6yGwDrl/m4oGzkdRJmL3V2gD
+Ve8f/G2EH/dsfIAiAZNaMsnLzWCrhU5P7rgYZ7Cjok74qVvXmk1UKHE822AoTQ5Lp1ZTjw+oH7K
BBlQOhJLaEI5rU7KtTvUELGkFApfVrNqjt9RG58KM9rAif3HNpi/78UiGeulDfdAUINLBsXuVHuJ
YaG86JEXagBc+ASuCgkOCR2HD5+reduu5LuM7bF+x0qBCsElp4y2WE/SF5+9MgP9Pi1DyoVBfkui
ElR4xcEx2FNzdYkaNTNq+VQkjfx7OJbt7lWLgDUTgn1lyghdtBdM9+tyYW9TpBl+Y7szue3ndlzv
l9cQIgBYhZ0428FtWBuH0g8mgYDQIr6XfeLd/413Cb6hyjV582lRkYvh+ACqDoBnMi9ai1Uiw+CW
lfRxJDLZsqOzreChNBEIgtB/o6X2uyoO2/ynlp6HTiwNgayjAJEdC7azyMXaKUF2hBK3u0dcjqRY
nuuTcmEOnoQJVo6XxiJ7ITHzjmwTfFZzvyJbZdTtzo8kfK9W5zVq7tcTOLaxIBnPaeotOzpvl120
tBL5ZX/cId/iBkrnptB8/Bwc846Kokg9rp7DfdQ0bapmKKmpAOvKOk2ofr4QdRUjxv2bx9Ac9TlD
TdDt79UySyC4LBX7MUQyYDBFgY3tTopvd2EXCT6Qzd/qsEWngCt9KCO3cGyzZu6CcXB++6vpRt5z
jZZtbxXKKsRCehYVCLCuP4g9Hqf7sqB7zujwReCXfWyiKF1s6eIdDi3ixhry0nPJdKJ8wklCjP/A
pFgp+8P65hzq+nagcL6DU7MwIWNJX6d/+s1Wll3I50/AsN1+q7P78bsGSQOMA1QNr1pYhqgem5sB
fVlqd4fRrEkLCyIv8LRyMybBZSUpb8li+dsbepiY+E/NW4ynL5Ba7BHgxPIaqfmlU1PjdIdvV5UV
i3/ZR1V13jxtHZ54stzp8+QAaxGKKM7Kf8oJ1vceNJOo6dSLnHpS2pR0paua+Y2D+Z7erIqzDe1U
KlDVjgKehOB1elT0lg1L8Kq0RGArY+E0emrXd374TsA3m94Mx1znC+lkdMNFKXd6aPErC7+ie7LQ
/XeUlIWWF0QtIPmhJRDwdMFWSItmW7pS1WLG39fF4EY7RiEf8ipIUyxdWPrbpSP/hLJG8F9TxHWx
/rpATFqg9UoEXW2x1lXyci0UKBk0Ndgfo53dh3incsMKaQ9qTJBVB47j4hj6X8yUESZwl2sGuV48
S7zFju1kRlHoHyktsnZkJ43jU5McdV7fLO0ZOLaPY6F4kLNX0WoXkrnCpK+vm67eR0RlDXY/GSwU
vdBqaXglruiJOmVD1fzvAcLcvtYSf2SrLssXor4ZgfoLwSs8FhyCQpoe9Gu98ws/zHegTiFjuqzZ
NG8mfgRg8Fe0SFwoIC+wmzb9Sxzne8xvF0xijCNurw5uVI46CsSAkervd3W9EGFFd9l4dM3pBgRD
jIoyNT+J7XtQWILzik89NgGfObnPDHyLuFPW97ezxx2GNwB+qqyrw2sX32VrhrvIUDu3wPdpgsSl
3GQP9UoUaKOt3biRkCQzZm4Mw/Hls4nFDYEcd6CoImbApFMxC1wKTzUioSuGYOpm/slO0qAiX0SK
g0XJy0HIbUnSTrPS8vrC2d/q/dMLKCuXWjuk7U9j1V6x0F5gtrnXyrQYiJDDKf7XjWPR9TKo5u9z
RhgDHvXvSWEFT6mLJpEpdyP0P4gjun13cxdhW7NIj00RsTdr0K5qRrfCvhOX62mY7hKJWXF28LUF
NLQQmF7X1xP31ft5xmTd08CbCZc8WUM+KawcpdtWI7GTVv+9NoiO+MYYVjaWTgtSZCx88TtONfTb
ng/RvQQYTpZgaL4QVT5fVAMo7GajI6eyQrs9wVB5bFal4W/UlEIFmJitEYI6tD3jX3WfwiA49kfl
36acKdgPYhNyciQWVAGec5giP9lT6gSRBqTXUwdXbCeTI+L9SwEcNh8ryMJKSmm+TJAwQo3ILJix
LMzzGlHI857W7mr/xMCzVQsMYw6G0diSCg5mcyHNSrSV6w/xnlNFl7csvPd7B6V5mhBbrOhzkR1z
/XDPNxrbrPgZbl/urIPnL2yJDKYSgr2ZZcmU3HLTP/8gABzLwFXoco+0Y2vRy8vFeLffsDTuvqMX
TEyxoSVTwEZChFALPQqUxCHhKSeG1XZQ9CK2bxznSDhGtwdSYrKfFs0rNQoYYpJFkoN9P6+k3ISy
mOHadQIIKbLHUIsG6Xz+CKKL1U0G01O96ZQlQR5404xX9NpZVoc2KTvwKdb9aqJRH+1E2zlXTvyz
zGggArGK6yX/uHzfMwZF+C3JNLyL7uooR3uj8/6C9G3LmAxaeXjPWgPEJDqr+1CvhmP6QMWoJ/Vd
D7D5SfCJlViDvGzRrqxMN6xLCRpffN+P0jrbpiRxwrGY/WLhjZdF8XgKHfk/DmpDmeZYgBFa1VTW
f821nF4V4DjsIETHaPthd949xqPoLbCGXEYvc3T2A0qdin+bgs3dQeaR6j6mweP6z5UFg7S1zcLP
Tmg+MSGBQ7c1naJWRc9supIHCRiElpZ2jmoowA3zP/Pismf6A9DsckpI4fmKyIoIgSP1SWrGyoGj
r0KGBfVLmU1isfguYnUIqHVOtOEceJHZ3AsLqqS2L/v6oKjq1BdoJ3KizLMBi5GgjMv7BJoi3W92
V72sSAKLX2b2q1YHsZ6K13YQzWgBUajl1xsliG4Y+CLp3ABJZQq1YKOrz2taoBUhpVWH2RAhKu9W
ki1iZCfHSCGqTetQqc6YVGRtzKHCVmv6pzuI3mFBCQcQ9wuvOR2yQVs875GHAeFhMcmLl1Kavqxf
T5MoAEmmh7+BR705I04LEyx6/z2QIXCuL5vtqqxc7cYq2Oy6tttAcCVFLDzVuuOHj+pxV62lQufB
quKaZNnop1BSYDLeyekuJs2Y/RutU3kP2RTCA5CNcfArnpwvsNbIWNwOj9GRj23UPpjZ/6lqSZXz
bciZ1p4D3J/KQZ0T2zp4b2bj73UbZdyHyHhYFdjr+Bpd9Bx51dK5djO+KWNotATWThR//QOfbo27
XY2eDQLe1D30rq/kKmrG8W7xtApTyDSg0hpx9n9lkvLtWK1rxPkTrKR65pUY+BZ2I/ERQcSJI/ic
Bc825f2rhWxyVkqEIDCWaVAZv2dTA6Hxj0UvLRNC/aRV7Vw/OAWKH+15C6STjQBcgBbHKv6f0d3+
98sCQ6E+UJetRgGRjX1Y3eJyKQQJcFOWdiYIX1X2zM2PoXLJEu7ZfIaElBmDO459dKpBkQ9DCL1V
vD8yX6kQqxGewWXOTc4RRR93j4huXzLxecG4V/b69TMczP0QBzkO0gGV1GZ+HXz94ssYXYl8Atv3
gpxFjXRh5gfsWiPtNN++vxLIuZt8AnCJQMkjR7J0HnaLdfgjvHIANdAvEpyv4exAI9DT8zZydE8Q
eY/2Uxhg+juHRigQlT4KS7f7p5wIUZzFXkXMESJ3JMzqk1STaCyJ4dmVd/HZ+Pq0E1N2W1RXWEc9
X7Ic7jEdONO77WEFKq/GDoNNJivqyEpFjS0cMmOGuMjOJ/2t5CGYXzy52jbIlO9R4YHvFH8vW77w
R5AKpi/bKwvhrl+1GtuQXx5P59iadNcHklgRUJhIasezbKEit/gBAyukCPtFUexKHTz23L1JfYV+
bjbzOZJGaJKvxwjs5p2ZL8JAEo7gjX8ycywGoXcX+NZe5vB0Ip5bZODE3HDytONSEm040EcgkEvU
JZHqHd5fNYieSHZcDsyugQBc/TUQfHK4AL77bPRPEiRLr45LXo1V8gpEn3EGtKRoYjm7NGnB6zVq
tE+EpKfWeSPfTVZ0MoP1C5I06HKT6izf3uIPlWdLTXjbFgocG3jV43us80b4ZhPylvEBIp4ynRim
koeW/psuyhSsGq+azjaf1oqTvMDMZRU2N4LRhiQTE1vmijenY+SnHWDjHA7XHPsmFMd24iqS82X/
rbaIid+yRW01ZakeECl2FctBZB3A0M2g5TljBoCKvFT6XN8klgbORTfuNtq+6xqrhLsb+s/REreQ
SqVWloJNteO1wZlUUd2vQwQ3R8hiqlJGG9eXyH/b090yxfz5qbmgru1Ro+tC2dcgj2ZTqc/WaTBM
awaov4boRs3oR7JWvGqt5nU0S2uPk6epsoW+zsm+983A6q10QlyK7RDQ0h+gFyT3kVr5Ssw8UpKy
7IGyt/spYQpPNcMWVhFmb69AqVgz2C30OrwAhTlj0GrPtWKGdcporpnmIC0Lfz8znfPnS6sruy4J
wY7Elksp5+n7JeC0JojR/eZ2CNtYf8thkcPd7vWjPEiETC6s0RzlYBONqBg5Cazgl52v+UjQRmXW
i2r74pytNmGqrxPsATgjNOv0+UqfbC/OBAMqBwZT/prTYRsg5UIdCz+lPNHRivw3q+khTkoF5nHj
RxZQtlhXgD1QeB+XyTLDLbrpWO6wiAH/NsQBaPvd+7yfoRdTZ7sf62N6sRTv1Xq+wZlKATlpwRkp
7TkidwrT0tKhYLilXuEPnMlonzjWTHZqsn3I1mNHM3kfYUdlxA4x0uXZZxG0f8rCQeA4wmEj8Sfq
MFcIiWk9XKB/JZVGwN0ls0YB9vYCeVctEKU5MSa2CA4icA9tDMMCe0Miz0Sc/3tnaCXhS97Zkcba
uUfvgX/HbuitKF7jtxvyONM56NhPAGJ4KETTuREm12dfnSQrExm5Iztko1wsWnbQkvQoXj8SSpG2
OphtEXqp70yIXbbvkDmBcIu4nS6daCBa9oWCDQGHd11DSzKVR9n28CP7YpTqmOP7qylFPc/iMWjg
Ugzj/fBbc8iob9oa5nz3I0dBhadfLodfGQHMEj47WrZ5MX9jNXG+vqQqMyfhPBtOvi98tiaRMVWS
C8almJVSUlUz55mSCinW2jo9dP0QtWbcsHx2jvl/drtGC0QVAwIeJDOrSZMyGhRbrrkJRiBf0wvr
1ItSvANNzlmZ/XaP5prbRWVxyvdYrRNsTC9xlZKwg55J9QnXfTvx1ZwR8EJcjwIWUaZoXUT/YvM1
6q70qUiEpCJL4pVcIM8eBTAPUzZzohovBUQkEWVm882p14wea+sPhIyLr1EHZjbyaxiZWlYUXYOg
+GWlxB/iBgoUdXaBTHRKe4rG+wMUBIY454o4SR4erFMwT5oc0/LosgIVi81e4x/LBMF/0CGyJdLv
a3W5DXMHCOsj67hcNvp7sTnvzP/VIhV43UbVW2TbCGpINbaaBoyzMu1jn7u6DGOXe43l8o2y2Ffw
zVo7FleCKL3K0DCF4SIukf3bgKOwzWvU+3c3zqK00U2MkhBcJlW80VgUIumnVfPgyO+RmTz8lUlB
lmYrAKul/8L6lsKM/AVGD7PAT/6sreajT2D3jxnoZw4erjw94szy09iq22YNei66Dcc7IcYclqLx
xcnaYp5v/M7J4gLC4WIQ/6JkIHM7QAi0cepIQTgYxdxWM8E9N7iYGa+GgMgp+UKoSsFiSdVQVAFY
/sCI/Qw3RzIOYfz3BzjeaL3upehe6bVvTjBvDu+/8Mly/5jxLwZQ3UYDrC98NGc0tWvUAbIqR3cg
t+20m9qSVlSDdTqXDHE4He2qJCKDmeA+gC1ntCntUfTZgVGo+gWuY3JPRcwhMiEB1Gu4jnZaXCzh
h7iQQKRJjHiArF91aO5vyXwI2XZ0G90lqgcPxvxmLulMESvMjW6ukKkqRN1Kbe663PjmkTeVdPhW
Nc/XtNjrXj+LanxwppdAKgDqvqbFT3puSgCPgUjKuX2SE7ADfTrE0QHGu4JiaE4yoaniq9bEs62I
qS0eEsOXr/lazYM/q2Hgh+TJuIs7JA6scs0BLGhaJumBfQy67d8lHSGSB4OZTTAngsex8wtPx7G3
rsuZ80aqube/fWffa8AwG9JERlnJI+01Ni6eXcR47vhCQP60L5jEfT5CMF7LsGdxxdiWcCYkQy5K
1+Fm/KF8CmVft3uMmvKmXxCIP25LMYxJ4Fu+3PZSPTB0bLh+vG3WBdT0jE3c98rz3/UaZE08Xr2/
7BP2lR7foW56SRTd5H6h0fy57ir7f1QqkYJYqLX5fE+15F1WkE3Gk8fvY6Jd6wGuMxDoKP6qAR6x
R9yCT66TuBT3wXrmWno+DDw3BqVBgk94fVtNpweHCVQ2sbbxcE/COy+O3SMldedDBBUiKSYprhnZ
rwugMsT8/VgQeZZZgaRZgDE6sj16teoq/Zhg4H/z3NllOIiXJ8YvhBRyhtl1wZHEqObA+HrsCneT
++tIHhGSN7KWXHcMYB2eXUE5vf+p8iIVl/nN5aVYfp7kXwGjGCcZLu0CLWQNuN2Hm2/89l6MOvZ+
Iff93FRS1Q6THwsqnGiFzM8ibNbWJDqjB/VSwwq7Pw8xIGSOi4KGB8XbeSGKx90l70KmnfG2+VQr
unVZCF51UDWlT+p+rp4CcI+cze5l0W0DtNjj0wjWQAEYAGQ0diDXkDW2auZ93FfJnwVHuPbMcDcu
S8p04If0Fz6b56z+l96NQoiQNOdA4QM1MwR+IkoOkSR9sEPy2KEnH/6JskaeUKJpf/O2tHde7p4z
Wdo+KOdTyU09aQ/vrcxWpZV3D7HB3r0Htd4y09hnH9LmEPZggg7Egq24WMRG5TLIH1Flw4zeI6NU
fMnjML/kehUrHiCmsKlcHwlxf8N9IoSAJmRBB3BWz2AZwPZ2vKaF400g0p7IZNDVl9/iIkSVt495
2kadthRMQyF6G9EBV4lULwukvM0DifjxT4k/MuCmL3T8RfJFLL0mKp82THWKjoZ0X6vHcR8gR/mP
zVj2szy3BwlkkNLBrn5it6/+7795MsozIIZhC+9g+UEW0FNOlWQ3skVbFhcWM1pTG8O83/Ruf5NV
5+w7HKtHiW4IOdsQisjX26BUqlBE4qsoOxT2TynRgMta02lZB9C+Q7crw6Urz0GxR8SmF0/+krf9
eE6oFzDXcg24jDz9yzZl94Fcn+d6DZ1VtXwFb5ijPz6rgbe9yn3PlnKPCBlUIe0ayl8eJAPIEutm
Jahnyv7x+ayA1U5/6BOaQ5k0c7NZuSLJCKsx8l+5ye2aqszz2FDOKdjfbMq4lHJN8q+2Nq/3xaPs
4u+PHyFIBAjHBGLCnh3CyxsxzIp9GY3wjcnU3pUS8tn8azqR9jA7kMvRozEngBwkcjpnA9T3rS1p
kzqPjABY7C6uwjNHR5+olbQX4qeto/wZ+Aot/fsakn0H5VgqKOiV3ECfWXrMP4oH8UVwUiwavhc6
Qj9xYfS7K9eejQpGZGOTLD2StvfdpP/cQdZ5BU08Cq5MQC36s75Pq1vX7K1ctbAbgXGWDSQ8+1It
yNwGdliexL2CFF0QrWRkLCFyyQ4VPXsjJd/itFEvOxCXOXcliPva2G981BsiMLtuw25Xr2EI9ULW
xXbX++iA8wFhCLWM2hnVzlZ+WQxyQ1Zh2vb1l63zJxhrofzF0m8nW96kdSAt2XLEwpPPw9nFwQsI
HhxV4GgpVffKy1xD2n6GUkx/oDz9w6DR/eeOKD+bAjcleHDBy7RO2ZzRL+R4K9He75XleF44Ubzy
xFICPho+U6vdNxDE5xgIQKejH7o/eQFHj3LD9qxhj4snfnoYBVO5ri6gmenAf8BSBWPN7W319P/o
XVqzuYUAPJOhh/ve4r5LFMV7N2akzNn4c81kWaj6Rl7YBgqf6NI65gHwxx9gsn7hWR9Noav5G0zn
5FxWf+ZMNdD59zzHFv+teix7e7fCDBwHlvhscJoEDFl+PsUGnsYAV9GaSLi6fBHZ56iYXKeQZy+s
GBdzOfadFcOCYGD/bb5TkKvM3RT3wYf9QppUCRZ/74mz34BWI/ow1ALoj1mWJ/mwLEPWd2HaJTRs
tAFX2/NfwbwWqdLjjlTjnf5xfdfwKRp3Iipm/9wGH6yjykqpBCKGuFmBOUJz16yhRE1VY1IVOPi3
9fkz5B+sxFI3FHGeF6g68B3HPpkmArJKliqlWlr/JBDmTXD1OesewjNgdFlXc1PGK6CWX+15C/2S
O4uAyK+VhNDBTkVwEq+6JgzwaK3qoDx5rogHKsrEDsDh8gj/XDPVNFCd6FYqYcss6teeaR0+UEha
70FnlrWpfVTdZfbW1os0QkLiI2FaSrdynESTCzUEECcXZzoOsP8520J22qKy8IK423gcpRPutlWJ
Q6cOFrm3ixX3iLbIWyMmdbT6mXzCdVPdabUtdKzLGrFikYRc3pnJ8w9zGdE53ihjbou2R9MLEx2T
r4O3s27S06QFzY2oKFUWIQJBF2q7TUbavFf/nC0jCTJCJrQIy56qy0XOz0+wH6EaeJQBes4xu10z
5KKGUBfxdEhM83Uu+BUccA8cHTqs4lPbjldp97UYP0B2M4d55mCf67YM+onBTXXf/b8gt4bbml+X
KUSYqSsARo/a+89AKK2NlBeSpw3XRbCosyUEfGS/den+dse0cFko4VPjeAJZ0wSdOY3nclxxMAre
5pxFZLS2N60IcF0y02JGqkHJrYlU/6vwYJE8b/QdVV/ITYtUxeDhBkK2ujYuwhG9UVgC9kmiWIRu
v3n/j9rwhpQN3jqa3/FLraSyDGBzTklhoWpVVEXGUWh8RkGF2+3tEsnrCN8/4BDEAcYjZ7aOXNgh
xytceijHsKjByjL9tA4J4S9uNCL8YM0aVB5IuXeTFroYvU4hcAlVXcf/cMYj6FqOiydvXFxzB50o
KATl/3F1De2lXOH720tZrfpKJWQvcpbdNAdI82E48nil8dpSLceu/GySVXGe5Oxpgy6SGT7hMXTx
eRF+i7DzUFILiWsETjXDWtsAozg+NeSKCJd7peBTMsokSenBmsa+iqYI5El6Zb8xSq6gIh6w/T9D
BadM9mOnpFkfQ0bhIepitrXyV++nAtH3RQ9o7r7gR6VxBPkwTMEZdUiQHIRZ9aTP2MFLWHBvZ0Ri
wYlmcjZBB4E+U6q75zZXZEiaZ4ax+pMA5dpgnMykAcqkD3xqKaEOU1CoAVyJ8pA2xxyrVt7gZVtc
yMmb/z5DPzwnfQg6ymmqQ6CKixY5oeENqFOufqo16f4dT4VQqpLXcML+pfIto7mmryIyIJD4VhxJ
kwbrDaV08zjXIIEGPab6Cpl78RD8I++KwdDIhNEGkv5rJxV1Br6I7IRa8qnu9fJT1QfXu/EoeQ32
5En+6UD09MwomZACfDYVehF2+RQLNoDvWMt346oSEO17UZRQxj3NIH5G4IjRuDiDdSoDNin2x2Xq
qvsn/qXgg+5M6N4dD1ehwI99YPUAgeykv1/m9hLnTwZKh2G6MnwkVXzaHC10smIHtdvPTeZ1kFx8
N7yyxqS43D+5pjXlM/0j/Tz1YVmOkrH+yuz8Rwm6kKbAz4m41zrbJu744uZzs+4lKoOBZxSonH9z
X0odNYGDt1lGYhRCLDm5hTFCOyC3d515/oylgs125U5pE+VIhtGddMRqNYOSSEYuTpaNf3q/JYlT
rjzNX2jRoPfj8LVLJgH5KTyOjvfnPbIUZJwmhFdG5yYZq4Wr60GZF3co/SccT0cfZhVdUp7uSmgr
0mSDsChxXgZKHXQ31tjxaHks6Oqas6yX6O5FjJ/Epq622ecXszEmN0nNcR1Brg/nPtAfW8Ih9O/t
ThKiSt+yUGbzvF2tCSiU66J38vzk+RaLyo96ctD6rES5bmtfAbduCqUzM51JeunPL0cyDkz8C3QP
HtLb1jtro2/SAWnd193DhVFL64r9DbUO8uuZjggIOXoDSA4hECJ80a5sp1wiMObAP36Du6Qeht1F
7Mk/0PQYm0udmB4jweTD693GHXCCbkhIbzEafQwv8bKbnYM3bKIYxa9OcPMt6ufX5Topb5MMFlmJ
qjbshofJihX9pCxECp/pNeW5C4fS0FOoYZCQap7TqmqRiCxcIrDogVayYQQxrV6/ePljZoXtMLkc
MgUcNWQnIuWXpso+g5ChNZO9I0IvycCg4lG5umXnTtK83Ri94ggv/lF6VT0lXVAk3vevcwrFaOH/
R1A6htJv9I0qnKB3zPP2z+A23VGVqE7B7zfeA+pgQBC640h62q7wN1xIy+Ai2icAwzCf/doOS/T/
Xy/qJEgWDhESmwwDuIQdyXUuBjtE2xllaviYR4ORB3fgFmpVjD77Us2wUJEzrkVBq4lvLjySjQCv
d7e57R14Y7XiwAU/7YnRwLMDo/oPMsc9SCesC52kZza0l9yIbjAmcb1OemRzR+b57qBF5v2AQBa6
tJCDLtPLi0Urm4iG9Q3zypiz76VwfJCahA/7mdiwc9p8g2DwAEjSgYKNffMTPkLIMgHrGGJVS43p
MVY1JZHiN6/jAzGolCg1ZgaA4MVBeIa9Aun5D8fIwZAwjlmoHrhW7g2SeQbZdjfApqR2ohAIJxfx
TDB9eO9G5/EE8xTzaBpKlvo10N2toVFaNdlJ7YJbU3yoNwwnry0l1kr8G0sh/iSf+EGuMB1EQNKi
Hf9QmSQxZf4a/dAtJiySxZ1UQ+rjwLEUFZR6BatWyXqHkdRmz3xZg3e5d9O6gFrhAFQuH2bgJrGv
4R9SqLe6hfl5dh0qoetq9cFNkxoeHPciqh6CFb861YSxHUyVzrw8g6gTagpWQe2GwszjMUNA8w3+
mVr+FO/twoN4B5hXlpBahQkufXu2te0NHMWJVwz5xs3opdwxK35AjYTxfb6DyeFoN1wx5HZHAzoR
R0CatEqbe7HBQ2GasKe7wm6/4aLcskEs/s+3cIhwZyaMjlH7f83bj01pBhu+vmSSrWOitpBUlK+5
wWiOfe5McPgbVd52loRgcOcP1XFqhsIt34G3qZB57QLexUeYKQ2TGmQt+W/GGkKz7TFdKYjXr9dZ
ZWzWbJz5Wg5JLpY8sbMvebbfJZxpA5lgFUneB4RCY8Fml6P9TX8xu6vbLEZ/tFj6sMkqnSYI5ykF
b+OjGtdOfmpGdOG5cyhJ+HbbcBcvWHb5IXm5lBFpc73iUsK+DmyuL1+VBK6azXuSsup19xsYEklT
PFGD+hZi2fhjp+mEiRrmqhY4N8pLF20XQ622zYewtXgyegeMbCz98mdbifVpNlyY6yKh1hGvkqWj
vBLHH7LVsonzkSa4IpMC+csNcty3+i6aHCHvh4kKntJD7B/Rl6fccrW1+7OHMgPEN/OmtdpbOq5v
SWh9yUDMhAa2qZ+ccD0FawhhcFIRwOGsdKGj9HO/FglVdmnzob9GyNn1U9Ui1992AaUYMwUnhts3
VTQ9dgGtH531+mjiySdBmiF/2BMDXErJD3g56pAagZJKBNiTnVfyn/6VLhxYhlQQfWKAZnj3squJ
+c0ylqvEcCHNfW1Bu5WROW9xPslHfAnmBsgI2aj7x4QAfCtBwn3g6HTfUp7M3PVQXneKctK42VQ9
mci4goC6pXBzjmRKnnSyrsdWiVp7p6pmoYKV3sjXyb7YD7319IjzNYo57t4N8Tt719THT39BPQUK
zbVQjVLDl/ZyLGgIXGQ4AlPRWoFX/NnQoKMfGw6gUxknQge3zuy4CyCqXi6xiAQ5CDtOIkTTtYyh
ziFw5Pr0H7yqmtekpmikFx2FxNF61Ho39TH73H6pMQ8wzsZvXGncC48ddpRPVwT+twhEaOY3XlCB
lXgdvfzBh6bMkT9bLZu87jXzLjUDfdpcQal+a+ZuMMcAEQa+nPCG0dJDVOit9n2j+GFZXy4NMOTe
yBtxiIq0PUXeXeluig2HMBiVFDmyuuFb3DbDM/7OgpJBZlYC3oB/y2ul+HUacU5eUtH52a2X66Bj
3o25WyOPEP7XvUFJ2qVMSPgwNemwHcJRX/52h7GFlHssXeKQyDjguXICiD9iq2GSXiVvUNtywwgY
LKxeZpop/AxhUhs6PHpdFaSDtR9j34WNSpImTPVCMeS45Oy1HOvZ/tutX0koV3m3ID337F3nNIC1
mn4j/tLT958hyuiOgKhVmVGuhI6pHgUT8jrJyyzlTBB8p4mL5iXnDUgBnAAxO8aJ8SPxheyxBuxg
TeUFq8QXOZKyfdQN6H7VUdHNU3bLxUWgGhDnBu9/zl5sz+fEi5HAB2Djt+21J0+vSNSwVO8X5/WT
2PNaQvMtyHYd7yrk5vqLXiYkeVybvHajhcmZTatH7moAq+A5G9pQlwI+x65p364+ttyuZ+I8uvQu
YOEdw22EyBVWN//5BnR6gYrDgdkvBjS1mOx5yURomqSNh5wex0f2KB53qcxNjT3THmvOgS4b2ZNG
ThcpZSFYjIBTOVtL9GzTgzOkXdvSdxSCf5oMMtOwhBZdlrCo9C5MhP+RIaA3QHrl3a9sLEWbNn7J
D0IYEENepLfZSdWPWlCK6gvbaUhKhA72RAY1n9PqZr6qsluY16aX2wgo/yIMI0Gik9uui3uVYYq3
WyyP9cL7Xf64OQu4GIO206aLQL9jwdt4lz8byk899qc2oceUgd0ENGN/WXDesnBX/PEBWg3XvPQ5
tptIy5fowSe+sCyVr8CJB5bFcCvfqlqLOzKZ7E9wq0U8bf5cJWa+frcK+tXmJvFg0Ys1z3XVwsij
3426dg+xaXU0PlVfJ7RbPlzRj2jd/5LQ7lW91GWIjCTMKYUt4hwJziZGgqHpk0mVUQ4ta8AyV5j5
yqxJwYvIYmV3xAUQiXUeLoGQpxL0ipYs4nbVP8luisToVwZO1rC3P8c3FSTQ5weviRcBOYwgMpiV
2xY/h3okbisqCemwBTcZ/WOMVua3y/raymcjIEph9QfCDp/aGWAi8Uo/cXZdZMKRMvolka5jxcqD
szVxGE90xi7OphihN8d6RVATQfQQaDshlUF2z2aW41gkf3vS9waB65sDp0r+CopYyEjQcYEQEJau
7pQgwp/8KyHBaonqAUoevCc/Nxgra4njBjS51aLiULNLdXMUvHRUleScFAMrqK2qwOWGPDxYX7xs
TEWcWXs8pmf3KDUXEksKGZNRxCj58IW0FI1bt2210it7oKYBISALJZ+GXJe6L0PD8b0kgJ88b/4m
M5vUObGm0HU+1lNhssvd0tzpy/Ry1wN+tTf5QodMvCIm+of8uGslX5ufiT1ow913dHTMCAmpAlj2
cryn25LLjjFHQi9wSsRGR/RGMsiui2C9qb4Okh9rfmvwFM2juAtC3qAA976HciUsZiEnEfuFRM6i
KPOQX2DUW+Es7VzFmMRd0lLnOCW08XW9Ao9brYpG64jFPgFs288AV4kS0xJ+jBTDd9p5lZqYwI+L
Nrhx+jaR2D826njFAoe3K/hDlUxA5ffgnSRLXjLQuD6JWngkdBrGycC5W7qfJ+yGmMXdHBmZa5nw
OjiJ2W/3pSdZfqHY23rjoE5NNIqumSMmjDmtbjssQEQuQrndeJK7PZbo/E4RVQ54BohY7ded6tf1
VIzl+iksd5cjAaSszMw0UUrS5daucIZt2CyzUJg7w6Ex+vGBDkHIq1fNyVsW5oScu2o7nbm1usAo
y8WjmcEec+2EaY+HYwLSu0rdA6uxd9DcnQ6R0Qx4AhZJKUsDg5hrz0eWd71LxnGX3MokFcs9/oS9
ZMXbZ395YG5p6Lpp4wZarcCbsmRfXqJyz7QjDGSsMyHr7z2xoRSSsCnbxOvZfrcnFdDiQM7fet6F
ZnfRaTkLbRCT1cnS6jUd4O68Ckn/17Z6UPG0zMNKWrvyP/RyL91l3W7quZ1gOu8HpYqYS8EKx6Yr
0V0Xjyl0gJpmho0qgoLAlBrmFc93Lf1cRGzc73+e1KxvzpGr+2gNBXrDoPbO6cTGpxvn74zdOxEW
o0oPmCIoYNRQHpBZP8QIWikvcYeP/xeidpXffETwuHDGvTvW9DEna0RXj1A9cuO2ALyk0kVHyqec
Xp9I/1XXEB5aZWq+8v1IMZJT9OFYkjdlSvyczdPk9qBBjIguxe6acz0BHqd9K33pSx0cAbU6k08U
ItKgG9WhRbwg6sHEt68dgcF4AnETD7FrFALna1bm9Tvlt3UUXkuR93sjx3ByzBU2Y/BORpqy5gRk
EZcJy0i7eS97jq/eh5fzkz32oQN+NchqlP99d1YV2f8ueoWplJzbpqsQLwKK5g5M48Iu6H2nRrH+
KGsVMDzR0B5gwTuD72uP8LqLjppSh0Tc25tcL1esbHeMGHo+/nJnAWEvFxlqyH0Lo9OZ0u3vbEut
GlSqRRGTIcu5UdwYbSUi8Qo8yebt0yymFRSLmvx0fVFrqaafDyHaiB9V/hcR8PEQN91zZaKAMcKr
eXv+g8WGXS48AruswJ5dgWXpw8jq7MipB9FpAESYUEpg6QtkPZ39ai0v8Zw9ZMIBJK20AwYqVvU5
m6GApyTLX+VeEvRxk+EOVdb5qw0NVYBct/taWsAU88P40M+46TT/k5q73Ab+plgpBJoP0nxucs8q
AsvCQHmudLnTQFMms88dXkXbgnyIZ8FwAznPLiTDlIzAW3d78slJ61VcQb0sTnCzcs8HlOV3Zb+B
LAyQQgVuhT2RG8cZT3WI6X/WbjJRN2EkIr5pJTSdFkn9dX1W7r8MGrDqOZFobxxGv2+O9xYCd/Nq
f0l+XWbTGjeB2h7EEV7nRq92IkswjWY2iZmmYxiV93JWkzek4N4bLU4NQUtV88mf0Vo5MKv4Pi3X
ngfY9jrfyB1zh0PBlZU9gqZ/BS3XiyByC7ngaNzCfS1B3la86DaNAxdLmbDNkcvHr2v29RzLmuQ0
AD3V2O+D7/Y1M/8eNaGCZVDf1IHuUzq2+K9l2g9A9tpiQA+aIxdJvQbUNAqfF7nbYv/9ueiSEefS
BVifpy45VuXyXwAcBZLQYeQM3eOwbyWxaU/AOlNY1XbcDMhvBMVLzSOlaWn1FSXqsTE5IXgx1Pct
iLpuP/4YNTVqF9wfFOwCuqFiy3wdBq36e3yA3qYPN2sxBUIgoEtVh+3qxob3nlkKo/9FIiEet7At
erODFU4NqDf9ve5fYBRMI/9PFJ2G0OCsC73L1p5KNIpy82L7QcyD+0VuIm7+mx6RIk2e7RQo5zQI
+OWfFujzIWuzTw/pR8NcYlzPb7SMapMnovOgU9JkJ9aFeY5KudafROf5TwX9Q5ohEKlS7KRVB1ki
ktxTdHKGETUIs+6k6gbxDFRU8MB+I1je7VE6HcT4/VJoQpPGdDXYWoyMoJMEKXGnic4SecsgVHlE
Apzv7r8b6YBsHoWk7Sm4h9qFvgASD4OJnIApoaryVqrPShR3hHVgbXVHSOUNHVuWDKSXRl7v17aR
6wQC2a8Iqxp3Lfr827kM76FC1IsI/8FKMbTuRmh4jiiUbcvU0eQ9YBQKDguMwYEzbCrvEfjRqNrb
7uhok8f7kxHkCbdx2nhxdot/BiUB0S/Ly1Ua1Frhw5f5YAvyDU1PW9xsdWaW9OSeQbXJ/ls278T/
G2s3xeUj6Wtz1LTAq/wl6f1jmdylLpEjAUc7vkqTntzxPBF8eif6f7xQhIntq7fut4a3NAuhbwTh
OigRDnKVW3OFsXrlF9Aw5RAbBiUG0ZzHy6epz9mOMfZKR7Htpuh1NhACA6a1uidCL/dETS/iNUQr
/yuoGkCHwMxDbne/Nf5SB4CY4jQrRXGcMLbNaJF0TEkrbygOmcX9y2CdTflKHgB4PkQ5S0E2MZzz
a3+0p/lGtd3SWytSTX4gt1OazLRfMoIkBkDj8HSzHu9wcc5s4HeixhEqh7tv8a8d2cwoC4t79mB0
8SXgOD48IhvpJOaUsBK9Xhy7Oo8Rw4gy0bf9tPVZRXQZoOBqRLWTrrf+XTJ6e/1l3YZi6bZAhTXn
zWoYn0aXI9eDEp4nPLpXTCYcUrsMv767tjuITUwIBHrHWS0jeWfNd0NqSjJx9RvpjX6X7RDOw6aQ
5ATnNStveBo6EvkADprH+OlVeczjY87nCBdCCefRbjKR0FY2lbFpR+pcJVoM9OgFUbsMNlw07gFQ
cVRHjRJ+5SECDMoAOYQsjHMWvnWtOzEA6D2AJVr3zIHvO6Y6Y//62LkdiT5zv3ZFEKw+3P4FQdWt
UwIsAEMJoOe4wQ4SwyqXVY3YxypzPxtMFxPLcp5evff4vE6ML9FFDcflI1o0Zk0nWeha0d5U0P4a
bj4koAEpZyhwYCTmX0vNczi04LPxBNSOsedVPlpAJn4d/J+vk5qWjcYhDHKewNhTk0rM1ET8C4dn
xCip42yVKIxyxBHjAlf4ueMFIDy95sTBis4bL/C6e8NC782F8BiisA1H1Up25mubGSHkA4zx2xzc
9Hvf69PB/N853nzcRvFQkvg9y1QpIXe88AbjU4FRNIXB5jCmR9eJH9gVM65s2cU0qQP86VdN6KyQ
/Pj/NMkzvgq4wG1TjgybT308tUB6d/UcRiUvGJY1SpmY7zGuJRQHep1T9GaqQmI+1N0rMYvh71V8
N1QoCXoyUK7ucoc2vz5ysjw/oiZxTWp2YvPpOPACxGxR+CJ1jkRQnCMXcLkJIXqK3G/Rpkz35PaV
diZFgsWTAoXJB8M2lkHneSMra/G4wAKHkB56TRuJNaToRE3Aq6ikEqcNWcwHbO4n8qHpbwN6EdPM
Ox0UKH3zLMiMhJTr5OkWixW4eGs93WwrSZZ5on+2TamQ7nyPb5MO8zeUd/BOT2Ku47gF85kgcalX
8+y19AF6oYaGKMDR1TtdU2/VkkHI2QMRqLPNzYjWo3gFD8gSJTHFRRklACNazCWjlpfVQGQ+hY7A
EOrh3Wk7RVxoN0p/R9mUwpUjyPgjVUiN+d0dRJCwYSwUWBSUukh7NL7TXcbKt/RFrXHaxgL08yGu
xHSzzP0RunfsLpv9LwBnG0Efv+VovX3RPkMxPoeHGGNun8bvpHZqXX23fvhQYrR6zHhD4mlZfJBc
1yko95LPLZaA2yDCaiAj1+EUks3X+XMRh9lIpwEBrxYycMn0fIatAMhI01JWUa2zsyfo4I2O0N2M
d9B+x9Pnx2j6aNP5Im5OTN31MOvQorTRflyoy+mEmmz8B2FRS/uaD6oB39+Mx+VXH/HRmE30t0wU
Utixy982VuUrjYhGhff5UtVLPMT/hoAPzRup6erwb4M4AYW2/EL6Nn3AypRpciUYipfx3P7aEOwZ
CG/0XexcKof6tBjr/PAPfNzRMVjyLXBTIAU6ZZoVNawncYm8MyhZNY5YP7isLLv2EBAsGj9RE2x+
E89Tb7b+q9pG3ma8T+DyWnLT3LoVZDRuNViw2mv7qmKSVqJ+fQkPOH66CbbCokVLY3qcbCSADrPL
kVlDGL0r4ohfJlvQSGOAYtqmPEJ7xbRgG3jRV5WK2knfmcVTT4pDwdrfVjfKTvHp2ld2BLBVRyvQ
PvIItG2mAvfVRNjYfE78JaNiVMZEn1dUXezoOXS8gwMraewRtaGA90rl+u/HlYuhpN++oqyiSLGR
/MMOMhW028IYvNHt1cUKf7Rok0burE87ZV0Qf3WTng4tBZXQlwJKbv/WYNvn6naeswk/Mn0OTcI1
VII5Gl2tsymcV7J4OhPxTp3eNbcY4EXbfaV9js2x1LSL8OotRxzEXCKRKgyYRrLOxQ2sWRF0WLK2
4cE2uNSK1gE4RT+xh92rqjNBVOjow45zoxJIOb8tM0kq6ka8Qa95SKUh/tQU0TKPQiUZ2PRUcTgT
qYArdlWVtpQNKWmI8vvRiyphTFbhARnms25MWXHhd0vxNdcltt9JDDwy6dwlcgqeZolBnU3onMby
2wLlt1vnRD/09O5/8QdG8Ml6Bc1LmzXq5p/iD29KhI/ksB86UajQ+jAcKLwH7LmT1ox6CLgR9yTv
km3R2uIHRA8NoFCai4yLTD1fMfKfTtzArkhlvS1bOcnfCmAWrsYUCENs/7h6ywyWaLoC21/ibxXp
0TQyJmFpSXobW6GGSHQbjCxTTIEUKlXfrh02eDGn1KV6Xzx8CAPp5Oy909LMsuLXnWATAiiBBYU8
8/tIFnqfIOZrTvgKmzp3dtmtKaejxnClDJFZDn0XNPS08X6zRginlnMBj5aQckpbHL1xNYcQK8yR
dDOWny0hkfwUQa+o7blHum3q0vXhQKAhbfVFITVZGA+XQRk39HtQV+lgJiFaplVujN/emEcou9Mw
B3EX+LGoMKojFUpo2Z9SeY+CHOBJdA3mCQwm3EVAhjIpVFda8v7fMX6tybB8fvzGCUMjBkDIH7/4
aSZpKRkAjnv+CIxONbmjDIFfEIwjAOiVFn5uwKegt37SmGQ0aoQwZMSQMRIzpLDD5zcoRR15O/yc
jVJ9QdbaUh9NXANJHSuscVGZxeSOMVv1k9LwyLriBusxKxRgmdn0WPuiGc1VFDzahjfQbIPTl8sX
9m+NCW4n/GpjwOkGiMMOxdiTna8exKu7hPOwWyB8HwS7oLSjSef2neCVWcMSRa+fqdhUSdECXQIX
jovo+BRcWsIK413C7Gk52GNqOe1zkExqLE2rEbK60efn7sSlLmzR/fNkaFWJAvwF034Pw7ays52u
IdOorFA0bcogWMaHxyYOsI1Gf7bMerYarqOcz2mki12pBW+vP1fjTYwJsnVoLD36TVWGmP/gWbYo
ebFBYCjPVod/dFlgQTWVB8nDtAJCMOzXj6FM0gNVy6CzENxamnBTT42gB5Ttd+GEXi6/6Nmuz6WY
Qn6Shl7ajcZlOwq5iIjqwVSGs8In3THduL4fQr3PsFh0BR38psUgKyUEJHftbeQBye6HZwHqjBQp
j+boCyl+fYI8xauif4s3NOwcRZUDIdOzT252ztJlrHyn/WkWAKuR27KsuCS7o1A5eVQFJAzFvKGC
4wdUqrc7Ql+25l+MCQEGW05APzIT5cBPphpkivl88SXoWoHBX2nZCVe3MDtvszy4Ix6TJm8libgt
eo7D4hgVyAnYUVTJkshIbrAWgbXx7RoU9OvRNmFXw2LYo3H94gvQSAoviu6d7EV7fPI20eRH0Q02
UKkXyKPp790XixhQyX8GL4TSV+pXjTbdO1j2djnTjuUuyW3qkRwGiqUr95TYCZDVXkQdnF/V5x/O
ZUy9fpyRJ/Ezm1rfK4ih78L7eW0F8yxOdZGxlgBxXamUhWR6yOn2ik7+lKK9ViznfM4trMX3DvBh
wGuopeeNQpcEPN+/wnojpDgy3q/q5DVV/WVLqbClQgROHjuEePryO5J3odKM93nTIWfGGiwX5cYM
viq2xIG9t0sUMmrWOSgEc/apehX+K8bhJcWZiebTt5C+7f8s+ANOhaiLG6epj/tCxeXEcyT+qvFJ
q/pHrRIKhybIT4OfDyLwmiqRT3gMgqxlIc++GPVdQ+eruocGu3+YTKwYw5mu3eA9/mNQJIrW17mV
j45OO1Z1mgom7fiHT8ZxwFRDPwzmsUs6DVjM0HLb1osbgTdyYUNip0rv8QxmFjhXdF2miILm00gR
cOBrs/mJdn+TRfZ8492UyZySld2PDcnGwDYzI1OJ0HMpJGsJ2gV1OstaO8OD5UZ+n2eMBBNF3E+m
ILXkF/t0NPmtPV3OPBsrE+KPSxSSzg1IUcI+vvZZYvcLM2BeXrIGfpeljx68U4zGEG43JscOTAAK
x6+ucs02iaCxDr3cPkuUS3UIFwfRAuAGHKRlkcCGAopw/d+60ICvrnfvD2UnbVLuQ0wpWuCOW4YG
P4rAXZmHLPdGdAspW7sCsdxyKM1n6wx6N//O5SmeyA8U7+C6vWf+XEqsqYsKk3lC0jC+6fN0Vyy8
Y94VEqUbrv6LWHiXIoQl5yT3Ekdsyu4V0XFzadjNyw0/CKgtvgoYQnm0cVB0X4EpcuL4nrq2xhjR
DIVZRH0/Ja8etr2vRNXv/EwgSLxbWk7oIYAJVOh2XPg4dQB+p+l59yLUnjL9it/mdiOb8De9iV/x
cXtweN91Enm9vRe2Xf5WSia8mMaXzqxFdVsJzrH0rSrj328jyxkY+mNPEs2y7S6kEotUup8KjBx5
QP3IyKobo8IAgOMnT60PNGbLq6AFmnxZfs1VLakvZIBDWq2M4wsl5ct4n/yzDdc2MV0yKcDgyijQ
CBOBohIxnfHxXHZ+A00AknipZFpSkBxrSp4fjJfLNUliwb5108Hnf/BmyCDCNNmdYJmldNNKvWyr
Phr4VEJBG2TbWyKmIGUuYRUlFltFmV69jOtDs1LV83pp/EcLLpVzny4/TvIIevD4sxv+7rnys4xq
bMt/I24rwG7vUhWmDQBnF0gze5ojcUFaD/P+Y64Yj67R0v7Ep7i1+kXsIzaIPOKgErUG4fTuhuWO
MfKiiz2IpOMgzgSVkAaRMacpmmMN8OuTesN5EBa1kgnty9xK/AAECQtiaYgffHhZuflwrcZF1mQD
U+NsIq3kAzpPmb1nEutCPu1tpZm1CsmN3aU24eiEfisi8P955oCJlVaT0ND8jN0ZRe2XeiAf3QtH
bIV4U8yYa1rk56bqMGM1vf9n/f6avGAvhHMAIkDHGSkUOivITjhZ3pzuzHzNeW9VGAGQ0JKbkYPW
kaWUqr/D3qGPc57//B4yPIYLujo2ZXknKgUVJARRhbg5Ef/UXeDQipwAX9yx0av7oQ4gl03H3PmJ
TASl9Bb4cvZq6joUrpog2UxN3tOV5Ky4OpWah5UDBokS84994CVudbV8KTipSODr2s+SAVGPFjfi
5AoFup2YMH9bWGy+2bJhnYeA3buEcDtkIhoF2CALkG+sia4ZNZjIqL/CONehFLeR8NO01WkbNAWV
4rzsdPLtNaCaIYZuETOWkZrwxPLNvqdsWlSENWwlnXGHznfUjkYJ5mnW9qKmYSHwiSHGKerJ5O31
wLiAwVHF4jcMAYh3yJ4taiMZbP/r5iMhQHqCBiJMc1TZ4Ki85rfkWJKPYvQdhxMWg0kVBBMhvPSv
p872kDKMabaCbz8UanIP0QiTAvHg4Xc8a1y/Qndk+MTZFynPJuisnzmicHG7IqqZVfvRoKHTGfGp
5L+Fn9ljuGtlHuPWCNNq+HoBsIHEot6rTe3KaQBZS/9l28Up4rjlfRyX7tukzZtUS0EbvgNIO8Fx
jnQuGH4EK2yFyys0QhYj/xU3blYKAiJ/o9y7wtS6knZT9sEh36knVnQfg6XaY3T+xRS0GqPCEn5A
oXy5EL0iL34ZuBO7qpv1UWEPHNZxAiq0Mpj8UNT7sCYUql8YNTPKzivwK4uxeq7sHbZmUMreXWlk
WQXZkraGQMxmwSJwvrgwEZtuGMqtRObsXbo2Ud/PGpALvBt46/GZVtX4ynd++QHQi5tOT6cn8gar
gHfmxGCHrmBWH5JBvSo2UP5CHjJts1qqWGCVLB0nCr6Lk5DXDFXA2KSHLNa7sB7KKxi/VvyrzjHu
nhYKsxWbqjdFL4cWGTjOus3g33PqAukhNbNCVLZ51cg7umj99MHhAHCcWjzNfbiNgIKiK6uun2Sl
Ac4/kgHYcSGhLwsRUNi0qnzsNGDg/v0k2CLcAVVJ91XMirvjiIlPC5bTq+TZxeld/91SqL4oj2yY
sAzOn0AGwKjL0daJG1rhinr0snK/QaAhrKqBWs3QJ9SngCHBtYQwawexybetgOZmNWSwWkqk4yLV
Pfa7nUKzUt6ut1JS8zkt4lgoad6NWg71TJlGLXYjcwHt5s6lEd2lNgIYwHlnhPFj+YfudzKPLOUR
0Nb5UThSzode7+WLkAh5q/ZCY5e+fBoxuuRlsNl6SioWURtrqWKIkYKKwyZwDnqT3L7sL3vjWqAz
6f0e8TW2uycPLr5KFFQUR+JECFOlKbh9Qu2V/3KuS2vbJVAw/lqDuokdoTWxoLxiiZa67ZL/jekh
oqZrBFLWrkQGAVAAa7WyCWNLMw5MG11/krbA5DpZ0/xxvs1U9jkdnOiIQaISrdPSUcAs89M/0Af5
wvU8Y9OK/f4HRZ4ldKziJp3WhYyOZLPuDmkd+qkPmm3/5h1szjPAxFXhMGXFaBJAsRWPvpKO78y6
CksQ+8/vdf7omRvBkwxuXiO0UJBP3KTHqGIjs2wxskOTItVYC3xWnQb9pwlbvWHxZHXp40VbtdO1
jxnf8lKX/v/RQQc1YOCLuYwA89iyyOB01UlCzlAePRbSgetwPUiELk89J5R8IGB4bb1puHdu0+in
g5LC/yW0pK0cUFDVBSg6lsxLoojDU35H38McunHmaIOLdEZvzQq9hGXHSgZ/vUHUub1mCyUYRXLl
RjbrBjMAulGnsT7A35RamKp6pqtc1ZdXXxHDYF3sqZ93rDU0MLuFxTiNjVlbPlI6umiMMNRPEPvN
1YCpQCL1RYajPbpUYqLN1h/MbYNblptMF45sD0yuGwnemaelogv3ZTsXt0pIQvppObECF7YW9zHo
VbpZP62MlSj+BM4EOe6z7MYupYi1oPVmcgd/AQRcuvmrvj0z7uG6hdMTKHTIgTXMjRDz3k1ZAXBn
H/6d4jLxTR5NlRWxL9d89uyJ+f1i8uU8Z4z0pRCxKp8Xxdb2BN/I5gLQaoZ+iF9BfTQqp1/Iv02N
VdR5KtL8k8Stm4pL0m7ZC7fNtykd0WIYdpjsUyjI2d5TD1TAG66pVE7CFmW2MWPNxZzZSe1X5Ulk
W4QrNrr1dtQwo1ZYw5hsrJqEpy3Sidaq2UWmkYQqrDQqiXLNDbvcTaaoy+rQpB/CXAkkaTitngBX
JsrqeP4ALBNXNfADddIWL9ICKhWdgOhbp3eXCvzqckkpqNB9t8Bh5CcPYxXbeHS8MUHiOfGuomCG
WaY3H092GeXOVyDiTQAB6eUffL6tvlusJd1oipu6JmiRdCE6SufU7n22Aw/Yie2QzK8KXgjliLd7
8aloUPW6sat/Ydg3HT3d/Hvi2VTmlmkOtZbhdiLVGLL8M954YOv7E4zh2TItue9Ru2sl727jYV4j
eW+CaMgTlN6+C/5pVxqtO3CANw9dZvDunZ6CeoEUcT+x5VkC067YLDXn7rfHqvKQ/MlX2Qj7kHkM
vnPjZ9eAnAMI1pIRvLsgtZw9OcdqxkDdDeuS0TTYOZnF8xyFB91lLqX0FyjFD3xMtlZFBxvvWaGN
v0ehA3GcHJxW6OrO+khRxSpXBqAiUqij8t9RlJp93WdkyGEHGfB/9kRW0P90AwOQxANqY+Yc6amG
czm7rybUbQa/mK/xPCruEPdyLTIiOxvzeN1g9LFFYv6HFxV9uabRe1xru1pZTafs+gaoXvI1XZ7i
VdsSTIjlfOzXqiJLcTLtNdVvUsoe9yYymRd3/PdLULmDaRrszXz4BkqOF5iewbgHpV2exBDodZLK
T3xHRESThr2ukpYMN3IJD1kyQO1IM6voxrcjasyH+WhOL7x/iNkUSIBNSj8ldWoWo+F0fvWC5A3E
SXLUrFUqP6fgpF4qT9c27wOIN/SCLJ/9di5iKAs2K1RTpzqISo6T67g15K9ZEj6tL26Zn7WERF5T
e8FUDNG7aFP+H6vwjNAhAowciHH1H5NMuhqzjXR6msikOi7405MHn9r2uv7CyB6Mf9Dfp6ndXGgi
I2T33G4h8B/BlmKDq4XVFTjZC/KIhGYu7OHcaYKPeFNFJWJ05C4LDs1c2KpBDgU3yqUbrCb/lUAx
ysU8THanfJ5QVSHvYXcHO0XTaYpC5cALYaQOMsrIvFy+qQg4j4SIoEFxPuZdGfUspXaqby5k5Enf
pk7nj97LMXqAKDSP0K5GssOGJxh6xuY2o1+XdusDOWFIntaPF6iz1qNcx2QLeWEjnD6FNIVvegFV
CNxa+Q4GclvJ4bcMhmJAmlOoo08w5dr6n5MhhxOG2LsDkPkRsA/JcBbsqcjiL2yuTDJL4SMTUv3M
vsSLFjR0e2T4fYFqN5Zxr4OOAJljiYcGp+5POkcWdwyQf0EXQLeKI8Un739RrvZEnev7Bv1/cGMW
ZR59A2QWfMSyp3dkeOUuhIYLWtT2tficqlKyfPcu0nLLhe3gNv7221qnAscFii/WEApfmNYRQ5Z1
bxZtPy7ocvUdOXbmKyz9LmZWOsXTorGi8QqeiShNaO4ksp0NcOH4zM35XrW16VYMe0D+dfJDxOTn
f+v5YGQD1Mvq+rMKsqzs1xSBYMUICqLxBKlAoQ4xcrV0EitZ9UtshcvJf9k7qlY7f81QhxTKr6bk
Y2mf+5Xuce7TtmChNHHWpT8QaK2+Kdsk+t5bzc4f1Pls2aayo7DUJfNBYfgSSn2zjWNvoDI9piw4
qbv4bZFInf6qP+kN+XGH+wRVPGedEYuJupzk3JyhjfbU28B1qBOZ3v7506GE+HAxbFrtttT7YzQo
y6LzdHDY5VHhaGzxaB84a8ZzJkXVhQ7rRZhcQ2AtDnhh4C/JfWrwAgL/9Ne02nBHc/jvD7BEjvUP
rZzKhQR6Nr62++S5yOHnMQaMNHaunMyHszMmx+qAEJO5Di2qF+79n/YN9fSiUgACfJr7DxGCkGWi
NVxWZsNfV25OdaledkYmY76hbtXB5I/xC9EhM4GY40PA7jD5tDKwEjd9vDgkiGsLOlECWbxw+L5a
Oc7wj5iL5sIz6xpachyQottjzzqxFmx8n5J6hPwQVeG0NC3Gte38xAAchARjnwN/Snr5S2xS/LVc
QZRr34r/PB+DDw8JxOp1vd3P9PJ2oy8WbR7LW6rfx5qEEktXAXbzRVueF76yLoIGmz4YAqImxloN
d+P+kCmcEqD0ianHbg2p13x9nBPtF9YXYqbBCqA3Rk3uWB/9U/Ef/owr8E0/PQDLrA4VLL5Yo2fz
0IC15GsjkstT2py+zXv687IFTc6/y+jJ5FvzDxwODjIdw3eVBA5Z5ixeM5fZQjMEFxe70MPi/v5w
/eZOdoZfbZO36Kay4uB13UyQ5ZNZyAcSHtb4OuWP3XcfXTnDhQdxv6DDkoPKY2tFWtOPFteLVze4
0q2ULNA+EHmadHL1Z4MbpjfQU3E9pKbZ7WDLpl3jD1QwaUMJ0wfIgEiP9bJKF4Iq+lSMHsnQpK7L
lYRsRR68MXn7SIwnxSqLkuB2198TGjVIPZwIP60Qh3gjCBQO4d7LzEjW2T4AcU3bZgijWBx8cDTE
J7HSdUAq9Zljr35zF2ujD2uMvWFUNz9i5TDOIoZ+b6EW6yWShF7VaozXqWH03aIyvbHDs/U39uhx
uvdHn2lgR/UFl7EnwWB+iaKzrD2H0DVSwYBXCOEO3jF9nUqWbQF6KsvCRFxyQqFUqjkeyTC4Y28C
bYvPZ89gIiAz/wBkdJREzp4Ba1U8KXEsgEhyHQvmtLMDIYgXsQO1fPDSZjxhrgH/pKkjRiZzb/iN
Zy1zMftn2/PCdWK/khdYbvP3+JywMyTSedYyGwbNgYpzkhw6L6AmZxB4NNrQCTXJI1o0Z+cEyJLp
huVAY8EJ9NbpsYJl4k1/ZSKow585UroD4vgJl+G6dG0mEy47gQ+C2o0ClrB1sDz8Iby7I12YC9H7
cpRfjiKwHB+Itpns/b8nQei9U/+f8Xw99QFm4vpVKyk4bnq9Hc09tWuRLSi39LsbS7iMKFcZogl0
Vi2TPE34dpJlfxWAm7GXUmlAXBhhpoEsFmuBNgGMCJoMVmnSz9cpgqmaW/IMfsv6BZEAtr7YzPdZ
PNMRSCsJsrOmLBT7fQepIxjno4s5zkw3cGhJmhyj0czcOPsRJdV6xAdfrwayutfv7quQW5ghKx0N
MzFMjD9TO4LZgq/rCkHN4/fn8AuMcJEpvja5AubI1aRUR0dtS85zLIvM2Wuum+pVcZSVih8JzdV6
EHhDmeXdmkr+rtvXSlm4e1iiYKZ5VE7hYQ5BDZ+3Y3nemi5plDxJjjaaBn4UWbHkSWEwFdhYLWp/
yMxKAub1AGj1ZjkmJbNi/43I8WAlG0ZUnwpaUEk/MdsQ73mz31yxPelhOreTjumaoB3EdVet4bw1
uDMMOK8hr3v+BGTo+DT+6ZZHLwiRMT/vABpRc/bkhTH14UnRL3hmM2Ajot6oD2GAs0IZoP00mVCH
f1ZB90e28xKF+3gXSX344qnBgd9wYn8Ub6eozLOhMA8uTeR0wuyH00ZubtUlfXiMfR2oZ5nEdTIJ
yS2UvUEEmyd4F+pnlFyvMNDDuPyL6w/xxV32FyKSE9gep9T+Hr+dlobUjNQhRjb0WWCWh7AiZ2Ip
lgQxEUK4yONmptmG0BVpq/zM8VFc1A/XGTumTXWH9xphkZi+Uj5vIlFmvBSlUnOHtAW/lt2bCNCM
YJAVwW//kbmwtyzOZTUGmC1B8b5KJN7bkAPxxxYYFntmVJp61iMy8Yki1f2YqTpZUEVQipZ/4qFs
8PgM8gXeFRpGizoaiGAhJUzJMBZq1Gsb53H+ba2grP34iDYrJ3AT1RB/1YGNrfFdMBViatHhgdg6
wPSLE8rXYNqmcPqf3UerTHSUq7QvObB1tJ/GAucm7JvKJenKIS1jMbE5tO+XJPbKuQHAUSeZOEZl
6pwcL2/aT9yRfCmFpkQ7CRQ9jLnuzzE+tvuPCYJSLlOysTowIbUM1WOrFJD66Z8OuAuSfAUw1KDM
T0rH6RSeiJfHoDxebUt2Z1phCLbeaTBff2XM7R8E9flnMwwQ2fuSw0lhcGT5u8DlZppMzHJUE7DD
lG4ALfURUshh3ztBefPpnU8YUKzH6YNwmpmu/mGO9V1cSzojQe49BRKUs6EiPlpdUOV3gOW4oGz2
gUGKNPc5JLaEFHzC9Ji/crLpFAIqD/gYpsnzFJtA7RWhEjAEdTtZ7rY7uw2paUPYwH5hXkPUFeb+
LhKKYFCkVgz0tBGlnChwQv2jQl+NO8kPAhQRdkhEcljSdkLUQs4SlxEVRMJ3KpanYZcrIiwup0Fe
sGUuyozE3j1G3HcRuhQeE+Kd1Y8oqXdfbLyhVeQXntsHjqvaZ3X98NjYETokcTaVanGGd0sUk9+b
noY3vpJy/a6xZ9i7zZxdz/VU/lldZoLB54WbTmKEpngtaT1hc9sN290xFnIvY0FbdCgQNYy1BXWv
ookbyR4dsgEharg4XhFWgEfG2YwRwSAjYM1PZJNawLGay259sP/ciRIDwK5Hx5SVYFJOnUyEnwEn
igVEv3XXObNHEZAvixwPD4rIQXzUtXYCIVnDZCSKuLSy+tDdJXuKFU+Ce6qs5o+5zcIspNt6dLGC
tNYIrg5K8ukOG527djDLDtrB4hvobfXrawFFkuyKYpnzYyz1TbLS/Zz6YkBvvilStGbmfHp+9+zp
F/xaVVu0kyNyB6S2VLRDq71Fa2hO8T9gsqDBrlgZJWTJH9fRXHaRWrF/h65ONXLPyBQeZYLZJmtz
zzZXm0JU94AtXHyNr4Z/MVIPllTs+QhMPfe5oyHz5NaadRJ192KDzjPcAXs73/SmW2JkQQSwxly3
R0WL928UFZUMPaQ5QblvLPJ/n8TO0auDwhasPujG/NyDtrlF5IvwKJCNT7bDWQe5+aiqXtSH4Ls1
t76xle3T6xdGxJNGkAkUUAS/mTKUfWzl3ehxI5pj9enLTPi8xGmCFopNRAUxGcSpEr1V+Ea7q+fm
OzezmjqgMFN9RfABYzbD+2Nv+cz+d8VmzsSJx9bRC3JDIOLk0ZRSjmzb1US/JOa8S9dUe2bvKOb0
fCOcy03+cvl56YcwDz2o3mFm9C4b4mAMPYvuEV8RVbrcZOH56t775b+SiLR5m/7ndSqAZ8SH+duF
A5OUGDxfcIosWcaa2LMe2MD73xnsZHRE2Xoxm3F0J9BPyXIX3TxkG5RwN4re2CusknmIVG6YQQCZ
YpHq5OW6R2MdxxYr+7g/7ybzYCrEld9WRlls79XNwkRIDP26QOrKLABoEr1hoKnW1ZjcS+iiEnlJ
ARrkhMfdPMiIozRv3NNwDXgywD7ig21nR1t+SyAchl+MssivrRo4rI4XwO6xxDTQYk+TwyNvQ3f2
hOVER9MdgEq2h0COs29zYO1GH0NZUZUpOo4HCpy07fHVa9PpCNCgGi+VxgaV5BGZW22Q9WuC3LoK
+aXHEfkmD71hhxWvBm700/O7l6Vd5OZfx+1S4y10/fnk9CRwEW3k4I44TbwvXQcFbeop+EzyTTOF
htrTpI9+FwUqOa6jed/hdqbEDrL2EMM2WhjbDx9WS5rFwPnECf5uwkR7UgdGmR5Q8LHKQBB3yAzF
uVrZgCfx9XEu3SEcKrUfWDyIUTuqLZ256yy5+W9A7T+Z3tXrDDjlE8h/W88nU5sRH8re8293eJES
8EnWRjIvXiMY3hy3z2BG7hEzyb8HA4DS4yGXlbqK8D4YPfEgjTIDvJyEZc3X5JXJPnWONhx4oI1i
evVn3EjxlLlxid1xWgAWU8D+dMCKUQIAmhB176H5vvocPWJZVe6gbp+UlRGFRHsWrjskUHRV94RC
KXS4pouzFbiNJizYZcYzbkH19yhhXll/YVq8apVQHuq/inpEbvn+1EgTbBwATMvtH1TdV6pWlNhy
vLV6AQlmwdfTBg+kbO+K3bKhnoBDY2kJK5x0bhcV1YAipoi4RtQoxUxuxxExjB6f6KckTf7PJhpm
G1yAwzXxwn1kwdKWufSbJOGqsUK/RfnI6J/ZJQKGxguEH38dfCF0AUEKaVcxt3fzR7amPqfrW+ju
isRUp+MHLgjJvNuFXfOt+G5oB64VAPs6p9qi0a+zadBiEsZWqXUMbNJyiSCU2ef0JpM9i4B3sIqv
GNDP3Om0l9C+DO1iYPYxGmisTAHXKebGXQm/6pI3qOtOCvepFVGo5inuvC1mzwtrKrh20O8Dd7M3
8fIuc/KMSMkdDfpHo3NNrneCxbjqfJ6x/I2/WvTkTgEephx+V+KdTS7gbKSiCUnfAWHDFD6YPeX+
TmsS59ZpI/kCOnv8AxI+adYL85Rgf6HPD23bSYh+V+t4h7sPRMkTvcruqlIRX97+xQD+aE/Yk9mo
Qp2UimNovq7hxhX7dnRWU9K5pmULNi/PhzrsgcjlN9LyBPoRLzMhVVah9+YV4PZCfFEXcjZ+jkNI
VDtHYpzatw9tdsxu72TLk1eY/hYxSLJqJDmN7ym4RMAi8bP4iuVCNFqjj2R2L7I3TFcMGO5B3PSC
KAMPcKDvLSxOMRnLH1oNye+7GQfch9y7ioM2zxrJJ5cUrn5xKHcLtcI1NoA7jzIOTPPtV6oOOlf+
b5DlkmE0YCaBZUSycDsg01ueXMOBCkJA4VfHViyDMGsZhP1ypl3KELg5EmSvS+cqGEAsBTyPVeXe
6teQqyxF3cGk85frcKFlEXKE1ksZPuKqKIH0t4Wll9cIrjekZvV5jQQPVYGBmGU3EU08dAeMCHdz
QkItUQUe5Cl2XJ2ZTskD5j5hzf+Kkl+zIY+WDHJCidQ0GXtazEEVXGuwV9kGJCTNOPopkhbMbOGI
JpvHmOzwyr+2xs5HNQbdfu0R26zsgddT/wlTZxlHk5ScZSkZa68nov6DChVdO7mnMj+M+wBgEGW0
DPGqw9IxD76/3O0PXIVhtmCBTtVAlUeiXR11eWB+j3o7xTjo/WeGcI7Ch7zLjCpoRFihiWuRrA/D
/llkgx+vyK3g3m2Nvr4avAJvYB7k1/DDpT+1xkjjl4DDUzXscFc2qPhW91qamVF5U0KumGabXi6P
ZyRHMedwkFfpT4KSUzSGdznME3Po0wJFrQqL6aZ6m9k+Bvwd9n1hlb3X/tofuBsVfWxUdpU/sQEw
6/MWebIZF2OpFsiQBPTH9LSGOJToG0+vJe1JhSY8gAzSN5x6ReUSuKVLbRb1vh01gvVhC/1JPg8f
hvJxCaJIkbBQcEpjGWT+Cbe/1/rwbf8L1MXNTJ38vomD701HLajt2gylL+L06YJhSGucDifnTWTV
o5HEt7lcohgoVp2uqq72cfDR2mg+nLxrxUuncQ6ZTyEJfrrkmkzayJbTiLINFAMiwxgNZE2ldFR3
xRgNdYuE3Hf3uY8/jUPFV+HaAiOR98EwYROY1CrFQNwqAkjgOOP5G6jaGJS+BaDxJHeJDvaa8Zh4
/6Eew6fYN+zBGM0pnpAFjlpH7U+uPmsJw5Xe3NnfaYFafHGMrPkDi8W2xV95ajeXNqrS0aJcWvCT
R+YAuSBO9tNFOq1YIXdKJGkE9Az38/c+9q3FIgsNC+j5dngZubYQQBbpOAqB0mlpwkrcGKvlLVf2
ck8BLzls8aUa0WLASJmKNmbOEl8EAJGgCK+AUVaGjJr/xQhbk07WrP/yY9rql0pZDIP3Gb1uqDIX
xGCzjOpVJ/r4oXCaLkYkEH96ez8ztx1HVBjOs4dB+aLnUArdATDQ/qoN+bS/26+IBqyBQpi9md1C
qqnyPP7mIMXGDAG4n69M9a6JLpzAYouAa4lObltxvzJ40lPzyI0qIzEWq5HN3RLJ7bPFBxkmifwI
pEawOYSGINukA7uWNUujzQ4FkwX7Kc8e4BSklPIkkcRnFmRGH8n/q4QJfIHk4JH3asI/MLy5ltPk
vUHIjRSEAxpoKQIKfSHE0TMsU/AsdkkYesPewrWwvc+OVUtrLswJ0UJsSpGJbL7IY0JwlQB+GmAc
3YbcL0thbtJWx7zUIHr45FfBWFaZT7Rgviygo6XCZtH2bX06LMaBo+osPLtvLLXFQ0QVZC8G0Nfk
+GY/ecPPlQjahHR9UPSJoPfpe+I1upOBQ5b83oUqd4FbVQLHtXMfD14XicsrJbmZJOvlyW/b50xo
yRSQYt3fH46IN/ezSVYossQsHcum7zsyoS/KNczAjkC5+2Pex9fVuaCA6QABU5pzNgdglr3N7E5a
7wuLDVywcUD0/Vz0mcMgY1XCT+O7jog0rcah3i8sMJdDlxy2ZdzW5jAu6VowZNnFhdEhCvBjtBA7
wIZm+cMv8wFsYJn5TLqArGwNNn4JH68ePG9NzWTvZ236DBJwUa2w3qcaDNItY4VMveOm9D72znjq
YNAZBfd4UkO74enC47OmSCoIvDx5JVAxvINQadhrx9n6GOoPmg41SqEcAfQkjP9ptRjJAtpdUo/P
MX+dRNNV6qlvuV0b+RyLcK+D+NG/XChr9hh2qsATb7il3qQmfTGAJpP9p0JfsYnzYPD3JJNLuEN2
rQgtfyoko/LpAnwq294Hrt96b+Z9d6tptdPSJkvLqUT9J1KpxHu4RKnk5GMwrGpjj9dVhFQDry+0
WfX6SWjNdRqbNDa8z46agiERPAIiCExBN/KV37PJ1OqS3MWraKM0ukMpIr6LpdfbOGN3d/bbW0bi
pSkAKhWVU6KHP7Nr7vU48orvP3/YXd5bxofrXssXYGCos9wdQq6NyfCQ7KfzVLDKNgozBiQ8ifcz
iGOu9qfHfvg32WDqmWrZzIG38p7cNYN0CbskI72sB1lG6b1LOtnqYDqX7OPwOwt8HGpwoSS8Cwlt
WjxuicRCcmTi7S6iE/BzZjjgH1CCcoVGPOtWkGKRWDyWHses897yNMZk1IchAJqL8yII8IcxRZG5
N0OdiAWGlSObx6+lsiLeBwrrlPO+DHIlzf9sG96lZbdbQBTByx5dtaS/2elTS6fBYKKVZRu6EkIv
g4TjefM+xB307fywAJ+dycdpdmr68ehn8omxVW5JqQpxQJo1Xn5dNRCOzHhkyX7JqJpaSkNHDEje
gH/+hWwwEm7MqFSvuuQ92NFNgqhwU6SRhtSo/IzSJkAXKlJ6ix23Bxjjb13g0lwl0we9RiiSOkaC
yDHZwGVSH99b8WYqC8yXNA8Ka/tWEQNWED/VfPnQk6U5h7BceRsa98xx1pVZNZ+zLC4QgpBfMHkw
kKnPNBV9sseLRX4xJBndS1oHlovOPuwVAghRNWFGfVQBLxDSpyXUFIphzNcGbYSatHpmfev6pfeY
es3wW8aQjjI1+q2kNRnuiFDKH6zSda7F1HIZ0yZ9KgAeDJLm7OCpGQgU5JfTZ12yTaMIA6y+Vtrd
hXuEf/ANroiF37UM+cCi78i34jLojtLFdyVgxwFe2J32GU86OwQSrJyFRG9aNm3qjHpwk0K+8+zE
1T8a3Q+6bqVtShMTNXQ9PzMmrsaAThh22vTI5ZRL9EkI4fcmxh6BFxTPgcY/LmlxfZCQ3ZK12Dbo
THWbWLy102rl8gR3uoZn4RcQPozOcC7tdxKPNP6bmYPBvZ6kqdwBnrkxqtg9a2eWDpdQgPAeeyAl
laPF2UkHxkPUGs+y2eNu46q24iRt9knq7TzLC+uPzhdGUflkPJ/2jHcOD8H/aq5NEQ/V8NZev8GI
6lJTuIffDVbc3hIBw9KnSu2VwuU4cOTyudzVTFsxjt2RvJZkuAChQMO5BWpjHt5sJSe1C6jT9PMV
hSDhBzY2iWQZ09T4VNV11CyNNZgTMDDNc+fpWEwRkxfe0sBsAB0JLEksrF8tHR74BogZTWv9KRXT
4PLEJjs6CjYgTmM6i8/Hsdo4+gfUdjWLfaF1qH/x++zRM/xLduXo6lBn15/yOoSmO5pLTmnvoOAV
THdgziJG4Lbao7CwSbeABqAHmbEZbvHOg/x1gk74rAH3+Mq7NVGSHFik0Pi1h5GXpq+MvfWhpzKA
3IcSMm16AXyj1/GSo3UZ1x6wHFbDa/dVCanZqft8z/GP33pEkklTwwKvdy6SE/0FUaI1Ox6v3HmT
vNq9IhuT0K2Lbj7tOFllomzU6NUkmqNtC9QjM5g+nVs99D8ZFrdphKe/QJtWhskkuT68kJqYz6ik
048z70giTWhZy7xzO6mJlkgnKKqsrQn74iEa8tk6EAX+CUWBf1EROdORJI7gQqsxkEAtTCESJZYE
EsQilaaPhdi2w6/qYANabDhOJYNfPvWwn34eZtLw0jFTf8HfUn4cP8HOuA8cW/YhDbk803lasCfX
LU1TI3r1jBPNopf1kU2oVGauZNiKrCLRHNkBxklXPnhiqmL+wCjpkvm8pWODff/1z8chvxIRnedv
cZ4JDdyDKzU6gwKZBal0cRtWtkc11X6vnZTMxQ6ihqBl+uH/bLQl5sEcbIxm/2smNgAw56dvAMGO
QZVxsvRmt+1KVTz3k5juMCQojeizWu5Q0DpIZay/RqNw1avYef0yW6Q87NSaXspNZXHc4s3hmTLk
mgi9vOhmge3bJu8J9CIs/zyeb3EwTuGkVkRV8AEzURCOEeGL1JBCjOzmMyyqIvCiQhD3DULDvefd
XU00Abm79Vcoeq6dHEfRuGxNlM6sKE+RbFSavKzbP9rfZ+/hD4fp+cM00kIwO/jbzCxMygL0znjg
cX5hyNuYWxjezmoFBAZASWhQrJxcd21YC8EUlvfuGo0HqdLjC4wcZgvVxxm1LuXl+k2QtBtpvD6S
BTGHhLAqyTpii8rPtX47W/6C//i1MLhnlcGRlSmfL4SbJvq92BdjRgN4KVGk/rl/ECicOLgyULnE
RRLDQYD9CispCc8WH/lx95p26xoKcR4kFwRGALeiI8e9MIe4mk5FuV1lbMGOilpiRQ2jA/DwGmnQ
Krl3oyOKkz1yL31DL1tV8a5PFkROw6ysQYb5Yst6Hg8rdS7XSm0W96mKbwn/+dbmvrzTaNlVINQN
AwQa4uB1lIz/gN+14x4EQ7ANPqchJDX9+KNHMB6RICpSMZubBTYwliZAqt2PPAHAZmVaz/G/jbH+
KkaNjr+CWuRgnJf8np0RvKjrduMP+MGYMF+fsAY49nZHdiet2u5m4rVF0p8HC8I2cEdFKmSK30HT
pX88N8hL6IX/jertbyVD35tDXFt+azWOGzBz2P7kRPnI1LgZ7o96ApwhgFdVFurcVH11qVSjG2Gl
4QNhs4huZcjncR8hXj0YckMQK3UV6bq+lwSjQAJYBdSrrobDK34zU9DePgiP5uMCh0TQ14h7TrtF
L2aEyoLYXB172g7LUzQkAWcgZ8WSxa/FiBXhQrlk7gJUIenU11M5oXPLqu6cybR/qvH1xzDhM1fM
5W/bLDPj9GEhgPhYp7xlTkF1CO4JhKgQdN9CJHIC43O9QCD1zmLT2Kdm5rlO5MmaSRvVjZHl36M/
WGmBkO8zsWiQ/fGJiyfa5E53euGZEUrs46hUINZ9cEZ053x297wufhj7rTcnRRMxLGNHqKDZaHw2
fQxOdJQz/6OqULILPL3Y6UyGWMKyJYPSlLa+2GBlWRrNKMAIG9h0wVoLuTjN3jRlMgE9WZY/i3B2
05kltwWxXW9IT4DJExsVlAifI4MWpXpnn30a2k5k9kNSD/9NJG/415v4h3YTNGyVs1Z4a3bbLiTW
135CeDPVJH5WYazPyEZB/8hfvcGpFJ8JHD6qnd5maqj9OfVRpyNBd4Q0G89gzpStAr5dyedNb1ax
8HLsjDMz0Vxclu16QBOok4B2JZvUSPb1VnurqNH+Wq0m803ik/DRo2Zbu2fw1C1WnZa8ZrSYaLhl
Z6yZMxN5mTbwtbzi64LmNoWTg1NL58xif9giqwUKuO/YVUb+oUeLxnPi+Pd7eZM+Oz9KiodW5jTx
Ko3wRhiZ8sICeGmZTuXlSZ7SHSQuPz7AaZsmC+HyomO3RTGGCYADJcoTAHTraJ57f2YatRUvtAjr
zyGY5GosVTDTBGTR5jjlZ5wKBpSgnonZE6/46cOwYkqqHIc8tuHQ4xV9jwEFaCQqB3XHFNooAo3f
bpvvYMKrkIcr3o/M7/AetzPP35YYoQDJ0EXst94VKQYTqqhsW4PpfesSIY9kSzl1unOsfjNLSOqH
4VMqrHYC9XCssHWsiyjixMQr9C/2QNzvyzB/Ee+q7sLR/LZ2fR2XVL0fZSA0kF68eMl0/NnhCqv5
45uKVdJlvzChkQEXP3yrT1aqwMZvi1G2SNdI5WzVfKpijFwwhpkztCClg9pBWdiIaTEs+DgzKb1R
qhVdb1lJSH1nRMLkEmSh2IhuICw7spfOBl1UWjR+KQwV23fa6ArbJRXz7m57O/4uYU6UxtqOvADB
MEm3yRCcjvZAw93Z/w9JWuPa904dq6odLtHc1avF8jIo76pnKfxTrGxNAsCBfM48sdHB/ulOhosV
LikSLrrfV7wO5lo5uyRWW7+Aazo41baRBP62J830DJGBIzvOHYHoNO3T1x2HqjIABa75L7GdI6Dx
c3t+1OMhwFYg0ZQ4MvKELsLsAUfFgi+iUwU+Kc+6EXBt/NqZ2vxuSDJthF+xx/9RlDv3nK9PYTgP
X2w1ipwn5BgSRFArWcuTrieWrmMKURvhbecoS7Q69VeygKEq1+q0QLsbGsabN3m0U8eQg+11icxY
ohlHx5ghTNyEljHSCS3YPPNdZzMVenqd6u2j31wY64IGuhmXVDlCOSV03NVOpb8GgD3qXa75547K
r/dmQDnlUIJHF5SNNWMR6NwMuw2e1Z/uyd+e1yQPmUXmFB4XKIwzyhLTAhHIQsz0EQHjmFqE5LqB
ePVpu1Lcj5ihjKhm0J1EMglxzIDMe8zkv0b0LpwdYErlIFRshKRMvb2Gq7BVZbHqWlfcTK1+eTYK
CPtpRkcV1aHcLTzIDCk4KhXDe5hEGDTZbFiXXcE+/kyFYeUqnGG02fsl1LpIcTTgpXRdWAx4Ha4f
ikrzXu+oLOVzHQ74MO3N1b2Z4c9ergJOYthm0dYj4BwEoxQLxiYWNfnhGvdQwK703aWGgwgEHwBF
QdjD2deXypuC1Egqbv/908BsGNsFdFqDaBMZxA4XX2/C0wP06X/8PZmLen2P9j/BYYubuOYS1Awb
S9kUf8Hu8MHNXCIEGKIt4IcS6K1dHb7TcwUGsOOd96s/R+3wfodWhDR8fMIpxuEfpSSOgl+QNBTz
bbAf7w1NKvFk6j9TTRB/UYcXWVAf+3vQpJ/M0ZloG8XL8e4CL9rVT6z7pp3rmJMxCU+mFDtZNy3D
uRR4uFtywMbqxHZkwzxCDhMKIT60UmDQMer1xCkdWj0rmpSCjkzTSxaQCGS90RlnQXAPcS5/j2ih
L/fJUZ7Y7epwnLmPAjnvymhs5iB0rDInYYtiQx4d5o4vppyekWS0cysZkCfYeJ4gNd30v+ktykKZ
uu5J3q7jOoBm0SHzn30Wu+m5VKKvAGVAutLFUUpXrmHILjLCOjm0ZtD40K04Bm7DJtxHZLnGv8pt
Q3FjAF2Uow6Qew502fckkw4XNIh0K4RxPt4gIhNWl7eZmviihAMM3DfrAz/bvBWE9qdfJPjs3vQq
Hj0s6K/4Mq+pBJHELfHMlVPuoug9GGd/m35yqFG4SKf2tMzN9UWl1OMiWNJAaj9SgE43Q1TBSIbp
kYJWRa2YNYPzMyEgXVz3x/1UPNPrRpnvqKbaGaNhKd72VkZZ02pAKvkUf5izRrDfuIkuR+kuCZUO
jTWXXWoNQ93JYnjTAnJp16xYCMp3nrzY3Yky2g6v0XeuesX1JgFvRFQckdt0ra9pT/+qnphTBcz0
ZqyVojU+0X6iNLFXi2KkNU/3hDlyO04O/qCoPtGTbZ8Jn82laZWZF2VRE3gmBjKEFKe5CoDqqFW6
J34GQ30h1MQ8jSbSHhkpoM+s3rAlIbaEvRBLAp0Z8AwoUfNhEAkAkHwxta7vVSjCpEUAwPWzGZik
2OjhtzAmbGVZKkQ6ZUSxQQjQO41yUpi6CpNX/WJa0H3IKQpLfAn6nXeMwZv9NZEmLjpLX6kHw5wy
q84dVD3wWeQfqmJ/8/pKqdCxLlD9RUkzQBUJ4slngfyYifl1Y79WXULeLqxl9HxHvATUojX2e9DF
FaOpcPnRLawPXI19wJS5cHtgkPeX4HYZj75oa2uvU0391zbV8c6eXJEKbWIGYgvPEqi+0Tfq6kdI
rv4GJdVM8XOZEH/CUD5Vm2ybrh7M5YCYmqDK4T3BO8oSqAZC7RI0MafcnYO0+4suq8GPGJ24/DYv
WeO13IwoOOgdei9z4LYwWvzTmMc3fhllHc5IzudRoECLVhuoQCe9zgDTNRA/+0WGXA3PqkXuMKlf
ttqypDTNlOvWDFPZzTsZu0EA6wkCiCI+iw3pzybzcMqVDBDpldrxl+x/Q8dd2QWB7ZK9e1QZWGwX
0c11yvzsVXZW8oRy83eFpGLYRra/qRtYBPChyfWqVoFX3+wQ4lrQzovVCWUFB3x4y1kgJdG/BA8h
mk02Gdj3RwXvq5RoZk37cUgRfCkxsbx3YGEjAMIzrybpBbkmxd6jQNRbDGwi6NE4gTDh1IBWGkch
9Rsq8UCCd/JKLmnZcI6RGIOfpoVDXq2hQsyzFMEwfLxNiXmT6CrDUnpz+pp2sB7Flpis6LiS4OkF
N+dZDq83FRaRorQR+CSpzyoYwcQ9N3kYubAdnyYo2Riype9DdXnx/CwyTGKYzVSeo5itTJRYTC3s
wnKb3Gq5bv6HG3R+x2JohrXI3xVURFvHNovApdikNSYvJleeZe8uNTDMB8EPiH1sbxa6GtTvX8JP
dAcfAB+dUb7S9PxBrepkofQ7I7rUAmUFydrBCsnAqgZSjLcisaIQ2MS2TJQ8XteYmVK0FfPRSvEP
rK07ffy/5y5q2W9NvlJB5CsZwa11CJK4PhqNTffFJeYo/Sj3Dh8TeU9xi8u1wp10BEVagYIyJYw9
nMFOJntgPYsYLS9gbCR+n3oZ9gdvJlXtDXF3uysP2HMlBm6jxiA9Ki7L0gdZUBotaXmkutDxe/om
cwDKEsFLHS+EPtvVD++hIv7XX7snl72BjWw2tGmsfdoiYKhW0Q9FdCQnjAdBSVHy7U1a5OABVZN0
HIcYI0cm2Bk9jzUWBW4Ln6Vw2ievv0fbTdMbFLzZc9d8ejNrh0vikbZzE6PrxFWBS2pe36KJ67Ka
01b54zl2o/HmJtmmgSIqgxYZFSOKjPsLnbfwqxkoghGU/p5fwKbd4QP0aZoh457DhqloTibEXZUp
nC8pDIWtcXUzD/Q7IS/J/ogGbOR08e+PPqKenUJfrs561GYD0I/fTAW9TwgGQ5I4IsnxpRLFDPKj
AHPp2BR2mv6LcyH0u/h/0otRE1FfZlv8NCBgOQwMwbFsSSVGNjE8+/NaVvDgtmBVYztx9GDvdCKV
v3hx4gtHTXqv2HlSgq+n+UACgeF24P94jDhx32BhJdXC7/d9lhb/DFBgBiJwhisA5sHfvxcHL29s
Ja+P8129wg8Q5Q5BYFwJn7ANrSB+usFFAq1d9tvO1wshosXwNO7QaqIRIUQ44K8mipQrYeVCAcEY
ZzURiOuD61V+sCHrJ2bPDfAj6SLGLdnpkb12eEII/7rWfGKUbSLzdtqezBSR60SsUzEQftADK6j3
vj6p1BJVMB4/Ay72q6DDS7fCpjkUa92x5EQ6T9YC6jJhmIqzAzfnv/DJ0ElNm4YsurjBQ3wkDko4
XywVLdhRP5an7dgbikX1YH+h55TuklnHuJqdrre+9ue0KAht9PfJcz0aUxsltlrSzB3IRNGTqtK+
0eFt7BzD+dFUbCWVnEEDqM1DMODcFHvDs0C5GMdcK3qrVbwI9rrnVNquaPA+Gk6GO5FRYIJNu7J6
O9PEYnUHf8BhOzT0jap97OGLsL0VfcONSGP9TzLvO0Eo/GPEYW+lvOa769WbQ7XQ10rvycfb/ffM
w92ibovdpq7VDlF92516102ox0Qvxf+2YI48u4VqDT5quPE6GaUuyXD0BP/6XsgCOuK3YUHfg+ME
h/Z+6j41mvJwCF+eFRcqgdAPO2CSUNXBjdn9srQxI+WF1d4RN4V8w94qBAG5t44XtCZidMWv65V6
ta3ChKrAEvV+skwnCuGaUoSou0eyTVvG+cpVqta1B8JNX43+a8NWcbd1BMZTc8a5EUq2DwGGHj8f
7fdrdVN3uBpdAr7IbrjofDX+3Nyvr3/aP9pxs6wplxvISpCna32AwUtmVlrj/qFXTmgIP1jl2A4X
PwdaN6PQ6PuwaXAnhyAxY9u/DGDSkzMAJ/pUZRNX7buxSoMgkFExKgVE4KD0LdO7e7NFbHBzb/tU
Lu6ZZIhaDjtuwip5K4fjj6pFJRlhzjk8WTJ4Z7suB4QZuqGbUu4a8mGC9HKKxji8F9l7LxH7Kunj
6UMVIrmDJ0rXoTG7BFgVVR1GT3vcdpL+u+ZYVFAmnYaX2Zw30QcT0q5sA0MB4/LaNrG1qnHCrTgu
EQWl59T6HYEhSE/GtfmlRCZFTAbj9hwdpg4+irjI1Yk67jtA2ChdnPmDVHbPvGDQYKe39MGsBz65
zCAM+LT3H9QRBd93upbbmcUBTkFjVj7f6WWo7bs1MAs7Dm9xbumOQ57pWzHSZerZJs+u7HHsPUvI
Uw8aYa9UghVsLHVOWcYKBBmUPfN8Z7SSsWUuqQUPsLZbbRSZDUHRjAyqf6Hd8bRyfe12JgJX2plG
jFQFnlCzBJXiWu+jAK+ZY9w+M+xuuoSqazlkunFM4OjCFvspKvUFzZ+nx8ZvgHqqQep11qA8e7Ha
upHAfewBC0CuOd9H1iKEfxeD1liJABBXwdO3tuZXJdQYfosX+JQXYvqjUGHFaASPLevd2eqCx8Rz
2IkyObZCOGKA5vNmelBP0oj61d1eBOKu4SWGHknBx1A4evPy5I61Z2UnT7Iy3tV1HMyDPs4KbeJw
HMYXv7H/CS4sp4RRkY3ombFj4fgsnlVnQkylNYzmogUHEM+TJ1LLyYJ7PPMK2oYWYMP8ddSPSdOk
wE8uONAHw7oVNHgJECKq2uaMnB5T3WkK8ugE9kWrlEA2noAvBOOb2zOxIDYBHdPlNVl8+moiBHdf
VaROseQ181Tc4w5xVBkMPrkykQ+vLY3uJR8Vb30UagkfkZWsdqpBWlRcMKr6xBGEYoEvIl3WOBxX
bSelLL+EnR+EXLbOI0PcPgcwbKdtWBgRCBFx8kvOeR+yx4EYljtJzMrgxnsHiLlf/prYaXeqZriT
mrfrXiacCVgYN+upUhRa1TJxABZczoz4afRCKVWiv3EymhAe6kWYFFx1mJW2/7/sfFBiIIL2TUfG
aPA9AbbrbEV7Y2+B4QI1ijGQOVHa1FSmokjzFk5m9/M/j3YKThc5tHRNg6eS5/mt3DZKJtcwuhnz
OhNSAXoZV//5Zo1sgEbN+TYWgG6kWgkyq7BNmE8/S12iWxQTWl0LbVtXMRDfUbp/pkHyfuaQsPQf
CrDpM8HinWJnsgIfrafo9mGRiOARaLGd1WvHVGf8JfCWVgHCadhWVzGFYEBAooj4tCGJjKoJU6L7
VCc88SsRC4U+mHrYWuxEGM6YNGjUFEIuV8w6Q78ljL+ssFI9UQwxKzy44VBWFDKQMtHARg+UWDEP
Nek2UhNZf/NblAK6qP1+vYskDVDjmt+krFAm7WGXrPwmNVlTRYW04iWiXKFxXdtg88n6wwd99EBT
e5GORz9d4MQWEnQy6tPW4JQReq6TJkraQe8QkrZO1t2LIqVI5bHNnVTyjdaSck9YrZ1Z6V1Ymsod
HbW76t+Kt49t+WkVxESjub34ca+3PRsi7iRgezR01Q6Hg3ziEKrM1PstN3G+cH8aEYD3Ygngu5GO
9wU8vAg/1tmN4f/7f5jkjG6RdrVkE/cGZ6Uv48SwvXdyVovgCcuyyj/i9Ll4CB8dehw7ZyvjfX7a
khqBaS3JGFzF1jPiSTlDo7iPKgn4Grptc9fwSB/xifVcLSGNW54Kxwuv4zabQEluJ82Be3JTvMx/
Jn47Q2BkzIl8jNGw/bTdwvdw0cvJAKI1C0FwhUtcVPNGAlO/cW131mHwVC5LUpb7M4g0nNpf5P16
VKMYnebkaS1r1BE9iOfP8wZVfbnOYvha6S0KbswhUAdP+1eWeYJIaPu0H+c0Y5y6SvdFngPVJEjG
WzREqQHHpfRyOfqnyZB39Ju/hLSd7Qoc43ss1slOZPib6Oatw472kclLmpY1hSCVorXe0o7uGRzz
CZFA1ZLDwzWcUUohSDttGvK8v2VZiUElyceJVbpSPCaPm9EZTXrVASW0ey2q3iTBZM/FjJYZT5wM
VLt8QbyD6lSMsrltthWFF4dOq0Yy3NAywumGdcxdMayVYccWZXLDUsFskM/WdhkhYZTvcvzEsvZj
dyIlgsTjILZq2G8h5q13BqLPbBf2EQM0lZ5ASjlVbt47CQinWDbm69UWkFSi+ihWFgAEH73pWrWf
fSx8OQnTvRjZ0+d7ZMZ66Horo2ZSqdiTH1LVnAqiTPBDfsnpOo5yw71TtJ+G88qYHetg8rVyAOs/
jPdedv30L5VQbxffMkM4EVJSSBRVByZPz6PH62uu9sZ8oXuL7a09MtDEtcfwPcSETKqS3pc+bZ3D
ZNCQRIM0shxf/PY0ot8EpmWRtieU3wOCOY/8kxc0chiPBGSxFPg5iHsM0aXy0EKGNmMh+5D0+r74
MxSWQyocghdzkW67oeYN4XFIm59rVX1Yuvx3t7Nmt1juppL51GGOfXmMg3jioKIQddQhIKOhJxry
VyZ5IsOawITRr+EHLlvKswKHw//X99T/cva0kio4xWpMFbz8DBEcjqfzp9Z6X8gpGBvRHIUQAL7z
VyEUm6vTuGVb2qgzEiDQfd2pNM0lGcgWdSP9y/mdqu9qTXDyqSzAcCuclndoMSRWhYdV/722KFCJ
Cw4YGqNjoZMCsI7B8P6bM0SzkYr22gBfAz/fxJplL0yEm34Tw9hHEf6qBuHv+rJy61QjVg/npAX+
jNO87Uhml2Y0lddsqUaOExqVwCq0EGJgfm9xzdvV4aoVtDSocyPwJfgH+Qgbenecus28MxwEYAqo
b+tUugkN3L76Z7DgxWYmgqkJVchg6FvL24gN53uWRnUoWKsw0okvWnppxhrBFj3UOidnsERyhJuD
peVjahjxNSHt0WqjcjMuvPK49gEHpTnKTETjx9uFHYdsYnvhrrEhL1cFm9c0ly3nmGyP7JqjmhIz
g0hpzideVafCLjxmrryr1fSbqZmRDuV+60JSJwoksbSNdWHWZ4m+vngRkjzdFl0HneH4d6UvV2gY
x1OttyPBLXsMQbJ8XwWtpNsygX7xk6+6KgOU+eLRTo/jJWqaRYfTQqcqVikbkSxmi5AIfuephhtu
ee0K82v8r/ft/wumx603RerRrUUX+d7v6UAP4oORm6KwekZUhmgf7frroUJJfM/OkkU7cJhOMkhb
NQX5Ma3WM2Xxywq0piGLzjsi1PI4v9y9w3NbP+NIWa+L5c85W23VDVCx+CKfVNU7vZ2j97TZHM7G
5ogPQw5+TCulOIx4oHcnX6IwgvV1ctsAnWQBUwt/tGOuHgVt3k1V4bNCPvHZ8MBkzTudtUOVSYlq
xLtbAKPwBHHOLXEYQLcuIoqdXblKzi1ZBSlk71i4S4fmeza8dx86JIG0Qg2gQLGmD63mxGL195Ax
6MIg08ym7qHLB8JYw4wUxPhAr/fbeTAAvThfrQsimkGs/6w+7IBGSo+dDCdJX/MtmDTYbGeS4gTV
rDHLAT3XRysFM5fb72zyMFa8IqC2QlYPvcSoADUcIlC0ZjpTWqh65e61epq0iVTIJfhj1AFkpUEC
4lY8mz2u2hLN62NNUM2dyBmvBQujJudgnC/hAvjo7vhCKB9JPOLbm7PXMkM0hXnZoLrKuFVAp7tG
aOh3JzEzX+tTixVFg+0ZEWve2dZxTytqAQdYFRuTkoefbx4GGpzwnMqXHEi+6d8H0yj1ZKztJPAs
tZuzCx3S9bnRoEV2dZ6rsutxjhZjsIb4LyWXNnloylX7vziX3YqYXW6Kj8RiAFDXsLFuocCo1Jmu
CW6xC0p0E1R0gZFiu+xgqhDOpXoOc7B9qbiJk70rGO48XCUWVVb7o0+3FJO6oT/FnXgmHSa2VWIG
Y9riKW9cScu9cBowPlh+aCbmx/RMUnSEgjcJo2MzOmMt6eCbhW6rNAhsXAEV3251FrQ22VgwuD8o
WYlNiPRjPAFm/2veypVreK8iAzFl0tE0Olmw9cSZtQJ2a53Gy0HfgrHhYM6qm2QPZFjyG/iJTudS
BaWRp8unH3u8q+oxt4HpkDOCwndDZteeuujw5Hck+R5OG6U88Vge5CeTQYguHRwwr57x4dnTNc87
CbxqC+z5EutM9E4vkQsbdEl4vnlY6juQM8xTpusu3XRpG0TZzqu4fsL8O2Ck1VIet1/T2qPAM3CI
rOOOXf66z2lFGt3sTtkm/a3n0s4k5X5Pwtvdqp8A/pyUhe73JlQNA+2y8Mio3jJ/82m11yPjTorX
KuN2o464uJvOGmOl3/CKM0ng4tEn7sLZU4pc1J1F6RtWc+CFB7Srubf/QMgbkha4HLlNs0KBxoSg
FXrlX2CaLufzwyUwWzebh4C/rlAFk797+fBHurwJL/5Nk4LgjgzDlawvphePKWWsKwPyjxHPiBAk
inm3NIvgjhXdtcAKasjjpTuf5wuYuSQX2JYP9WGdsy29PXdcVeuSTW7TKeW6N2Z/dixgYouyeXO2
Hvvpw2sSU1Su4YwO2fUQG6p2fo16cU3gt2QeWFLQZAPUXQ2CWQeJ7r8PQk4nKSTHM77NKG/CTa6N
7fJMtVEbS16r+P6uGCYzhTw5th6ZjgNmBGrM3fV6sBeZf9r41YY4goZwc74St88i8jutEZ34UGap
cIHz/sDQy4eZ+h7snG5TUYXlK03/a/IPNezTCOhvXPOchXnKRDGe4heG9ZZJ1K71EQ6Fso3aTvkB
rfcAPjXQ/wAkM9AmTtvewGsXRA3mJP46HRZ+mG07nGI/qtUMYeAb2zfnzO9UQ6XzMe7IgVAbHts5
vUojagFvhT4cIrm4lxscuAvvvleckYZ/1cUKrK1Co7MDv22RXIWEeEC7c0vXwIpCAP8S2BNLfzLH
tNFO6HYShlkIlaswWEiCD/8y1lJRTCl/R/iItlnqthsoPAq8IPZgso8DPbnCOI6BJpQ9ndvAMkI0
mNwyz6MzBtt+ctdJq0TqaCpmGfHgStvZ8K/TzjTGztYmXhyHi8cT7w+WGJVdMZTSUpH2NjMu3hf7
fqtIknTA0R8LtLyX8/WEgjN9JUKHwCABDONQGAlxeKLxvwLa5XBsQIOIzZNDv5ofl9z4JEfjm/lo
CjmNlYrj2YS7jMkVCyLh9BIe5iUMMS++sZ7OS3PUzXWNjFWfmOHNqaWo4UFYhMCXSRCUkKUIZY9z
HIiXvkAvr23rtNihBiWSJ0wzqHsC4sOFvRXugxqQKp9n/AicdGL3Svcm6PQQxvt3ugk4/BV+Z3hq
htGvLAe7fDrGfXKqv8TXDYZQcywb51NWjR+7m8ck6fHBJ4g+MHA9VDRqtwnenVYtHzYJbZi+B+GQ
rOvQ1YxWVzQ6tXTjEEDC2GawSIHsK2WiSD32+wazAkveAyrnBDgI6c/gZac22gZF0pNmSwGQm2v1
/LMDDlFPs0U90kmpsf6D3EAVLx6bIGGa0Z5cv4rRnmXHy4kWihIQk6Si/4JD7ENyUXkGY/OnubiA
qs6YdWoib1+NLnFs/Aa+eZIPGgPgloizuV95rg6prq4EkwjHAfZhjlkB5yBFM3g9bQIZ2tjcqCmV
x5uimwR7R/bJdmDLy/EDE60+mRKkRFX/bNkTJliLma+z0V140U9faiIL+6wQdVGhYa1LPgoEjRV0
zD9OPjDeEjqZRRo/Ov2Ziu6wwlo0uj/TKga+6+DOCAcgxDrXAGhAgbDBItBpg9w0IQnDZ0VCZjJE
d/QQC3GQjylY3SwCIo30cUrv/KaPG9VOISB2Quli7XlpzaJTlhtRTVtIH+7TPSQdT/PMvZ7pUt+r
grDnl0IhUt6Ly7gZW/IE8A3/M6CzjT2OsKxMwytkXlzbp+7ahH7C5tpHvpVxnlJbKYmXzwRDNyG9
Dj8gRcoVtXHnrO+Gvb8fBAqos5uRej1UpBp/w7SWzo8OlsX0xFV3Dim2q/dcNE+dh6ASdGls6bPs
aGPEcmi+4P4rH46USn2nvSNF8UgK4+3ucTFvv1fbycjAS9WSN08MCsNTbWySr965i11eAlADtO52
Dt7TCyggkCyvopujk60qjNDqSEUwZBTXsbjcPODxNaoMHisLqlLk0/BxLmOnxZGNM6q9BWUWhO2r
L8f/lggezQVmAZELE+yP+gqWml0IgDOrM8oIqEHybz0tekrDZjBS19YCSbst83H8DLRKL1TI0ceA
P07JtQpQDn5KXy/EypBxaoo8arjbq76VX+CjvkY1hJ2CVUqtGl09iIgOULLbCYHwxxpHa9WuvawT
CajA1GrPCIyiiC0+uC8vQWXZeal4y4IPZ3mXfQrkYK5iZO1aQ/emdNUJOD1KsDFBjEpTvoMMra92
nowJMXvDX2U/bJG/kN/oXTsuinv+ghPdfBrOaVEJ8zH3gv9pNzmFSB2yn7Lp82jjzjmQg9m4MNBA
8ZyJkbgSNjONwEKb17veJPVBcpM+jnZ28xdfSCCGN9gph5xGk9AH32OxiEZ7PtpORpkSAnbhxzQx
sFte0A9HAfHMtFrsbFxJKXtex2Pyw7o0tr0WXdSsnkSHkvnqjom8l8aOkgxlmwJ/Wv3/eUGHGAZs
+TRnb9mjJMHo4bKxx0JLXmdNb81pyb1ujzW5lVm9xbPWJ21OGLkd4ea4JMx9rjIbXlvleR9znOP+
JQHIpRB1KBeMIBhp+gKBN5gm9Q60VjePtPQURJWo++B6S2EEafR5rgebfqvtD3dNNG+C1raF29dD
RuV43OitCQt5XBeuOKBSPpd0zzpwTPURCcFTX/1M3PoslS9rzN2kXPXcCU68rCiVmdgbx0MCrQKs
18gxadZBcm9vmli1/xfrJzme505tm+MmDpLSGP7jiQKUP08k+Ey3/ZCg4mGomS5hVwhUCMd4biIU
hr93gufSmAtGWd/Wh28ODVknBa2LHmvT2lDVHkQUxZ99TpCzLJu7/4gQS1PcNEYAF6DU6y12jIQ/
RyeFBDeUtuDBFL00UTZglYH1Fx13Y70qnPfO0hXFxGGJJ7Z1Vdaa23Ui5EIv54vA94KHStRRt4Z7
p4RHFxPUpDgqLZYehyCGJ4E+3ZNZxYibPEhcc9xSpi7Hf06HJtjM5Osozj79W5OmKm5yYhxTb6dg
vxmgLEUwxwOBxM53qAOrkQT/CT30tmbIBTlfkzhnQ5BXR/35kNzDWO0Ja0aa1HN3o4loDEYyK2el
VWRH3nTg0kvpO7F2B3x6icoBBxFGqoMUt9QBj/KJtje82fAfkja2i1asHkUfC0XUp44d7h8SPy7s
0jaW5ZhK3jBOKqzonRFdRuBKeFZbcv4kYTAUHj4Jf09bL94JeyzLOoiKRgNKJlOU97xWqptGUhjX
9XV2UcHfOKusHpNb9p+n4cD7UCG5AaL5jE1J1dYqcd4Ih+o6mFCMlFDRq8lSAyXEdhEkRVx449tZ
EEY4IQnfZnhVsucn8XCopZ59ePGY9msJPRkEkHadMGb2dasUKilmdnjlgpON+VegxyCCeQHAOfnp
X7FGdJ1rMf3MjRP+gdaEbmwl5LnL0ig9jGNLwhB/mEXVmkiw7arTU4ZmeAGIO75XTotOZtIYagwr
qLaoFgBF9XgHeyVeVnermxsYUZqooIODP7xw/akbFxMZIKrjJyrBTStQ70g9uNv+Fdp3khve08kU
OwuKAWcfUmZOzLm/zFfQ8/Lo3Pv7rpUURYYd7gZzqTPzvylF6kFbO83eUxIfUWNE+N9h/kQwvsUg
xuwEkgBeiR5NPSY/6vtFWAftnPa5pIVD0dJ7K2X4xLzWkr6LNLF47YR8rPVwoa/4ILLqL5kxgPeq
OSu5eml/whRvZmdg7czZf/oeHZASt4Z6lR+E+C4jPRaxuKpVfDTsqS2a0D1yg4un9JIv4hLiSznj
b1JjYgh6zFNg/5cJGQJxVVNICegVVKmBb150GMZXrdQozu+ZLgjGscAHkN3QNkXRcx7BPoqkGjgk
tMX1yMsCEjqNI1nEkicmLl20Bppg+z13dBGJlAOMY/HRqW6wMFmh2RLE497xyvRXMP4RYdWhOsdb
SScwYTCncJ/jrxA2EuvS/lV+C94GByCvXwQKPuTjUjOV46pFQ9xuEH0+4xpf7syX2DmrrDeskeX2
dNiTe7k3uUvWc/RFXzVO5j1x+R2cMNH1nCNiEwZtpv9Be6qurP2r/MmSL2EMMdNSFsfz3AJX4nSC
+PzMnUkqfHxeKmaK7IVpwyl2+S727xVJhdnDouNuSHW/OGIGHu34tHo5U1uxWTgwMCFljYy2Yw7J
9gaY55/FSSyM0i8V3sYRE8Froonyx8Ba76Tlon2vtT+mFXRSgitYTuc5uWda7njU/ohPweiV03Sh
jYK5orCfKapW1h2QrZfU/4z+x/1wmbfwstqsKJk4MU15o2z22E7uNDM9iBiXAO6wPHanBJkUEdTT
/F2lrvze41u3q0hx+c7OQPgoO4DLRw+qDaja9CU1yX1JENEwqzzJH9rpPaYCIbb/H3Nojsv+P96V
JY3km7DUngHtpTaA6tOxUo0J8qYKAapYqgSOQu9L3uUpG4z7r0EFFFwH2GbZWIUAhECg7YkRhDYA
1iYNIk7yB4IlqFg4ykmebPh4ekPC6wIsOe5svrZt99QKrsNLm8FqU5X6jVdjV29y/koPi8Qd19fj
kRwiE4/IKoBzO3vfmHQ23fpU+doPUEZwnI8YkVdFcuX+ZatTcsd6OKjFgbKxCdz/IxG13WIZPMvA
fJtRi4SvJhPXLw65QOV2myKqPr7szEmZQwKrMktuOOgWcVRiQk7bwznVV00CWIuBKJ/eg6CLKnLH
Wxxo8ayranyMKw3SGARH+57VkNqPotYWrnx5Uv8GLBSrAd0vub0B0xGpAmLjM45JYL4pMnVQ/0zB
dMh0d6iD0v4GIuk9yX0r4Jyjc5pzb6LvrjzF7somUTmt+vtf3S7g9Gd1XkShjY0XJn4Sg49UZX/P
V5vdTUdvsvdlqhjVfw/dqV4APhVafH2qBj1mVUBAUFBYXnDSBsI6tFWA5XGdiwFuHmoHkgB06NHj
MhisoYv4JPVYM1T5FZYM1M5YAVR5mMZGnEj6wDFtc3bIf2ual9mPn7rXR4H9LcWRSJnCUZuXxqNW
xfb+HtPfK4Vfsb87+bOErp/hMDDXqgkdknAMf+bo+rXheI9fdCsq4sb60nVbnpLAPd/HaT+WOCyr
Bgo/+RN4QfPNHJr64SfHfIh3dzV4eIlNQYwewbpkL+60bBinGU5MpEQlnVPjUKW5/QXbUOz3oLBl
fGHeUCIAEhjEfCekSGY4NfUOcnnsM6DeIfcZXsH7u8ttUmtK+LMgPN5woXzYQByYUi1eJ9SSplYC
Nv3cO77ldIcTCJv0ezpqPqRv9R7QYEQT9cQUHcM6k+/FX4HmwoJFzcasBnuNeii000i3QN4bTd/g
mWlC9DMC97GrnltzsIpEf+9fN2kYNzVwYF3MrqJFEOqFYNc69+XIQygRpHI+Wc/i+tj2dDthBXbO
VtDQAuXYxtc/pLbqc9Ztx6roYK6+pJBmLvU1VdXM6/0wJ7SlDL/F+6mPBD3jaNYetbRoHyXTApz9
anHxk4PI5Q7tu3feL43N4HQQnGZ0b4zC+VS8ttTKOXDGpHH+Z11meg50EyN19lOsrRKMhcbBiehj
lLGi7Nz918/NpHS+XSq/pf3PUMRSeVyzmGyN4L79BYEs+BXZy1SEb6sQ3LEQtmEB2y9JYuWctE00
MOmYs4eUPehZzur4GuljLw93Ux/nNj5ysFisVbyrcIrPgH6tSQSr/rrheTXaJvQGDBj1PRVNHIr9
96lulNx1x0/jFj1pV05wpyn8Ljxo+EH+xAN1sxEISIsInbTgCsbaPk/w9kDVSfvCw+j4gIBoxfmu
y3i1x17shs1VSQyB9j0MNBLU1ayZBHNJVntp76pGc4DSevnqcpnedWkLuZ0mJUz1Etf8Md9rbKrS
owNc2kcGbe3qrx4wwmds/mr07KLth/XmIx5gqBoOREwzN8L1vGe4goy+rBpm/R+8++2r0HI97BDN
8uYR3Z5lui7aB8LBtMDfA4iYoyoVLFmLZAmJ9nbh3IF3QkKGqt7hRW/LarlaCGBrw5z4KpNUSXt8
cTMN9dUZnhoumrpJyYm9s3xBCJ7lK0ueqBrYiibRkT8+nkiUNA2c72wuDEikQMx+umWEzDlhyx0q
YkDMaiL2OwUru3NseUfJkuyLtfrs+8end3/sqVGYtFe9jmAh4nrE2s2qCsg64Teyn7KHZhnIwB6F
YWW4P+XUZmGLLuKsWjZH9/20tcp4vQquIu0RaBMM1fEhu9fRQr2q8uUDGpA3udHM+xZj7scVYjvh
+cjtnEsOSlo2TV/GgVhM4enWFrYcCObamSLy43icjoMegX/AIQfJrWaRlbQZcynWbEJf76sRra/A
QGtjfMZpKrotSklPQhRq1B0XQcezcfNRWGARA2d62n4lRKuYF6lnbfr7HlCb+MLugd8Tv+NqEilu
DsAQY9g0SlDVn/ri13KczgPpfbUn9vGWuDnVUaxbZdvMAg0bi1V+rx4zqObyl+lnaciqVYqdjeQK
Na48h8L4zxuBrtnIfvX8Yus/jbVbqlThsTpmxTnGGzcvzETnSHbQm9+CodcDaU/lpZYKy89xK6XF
vbTkxiaGr0tzbs2ofg93e3O+LaT/wwLpmgqWY2wiW80eeBgB+eiUuVvETNBmb4CWH66/3wygAAuH
K59qEtUJg5W8bahyHotqm7uItA832bznRRSE7JY2+1a7R6X5GlGRaw4kbbbofFlJmjpOCtf6BYZN
oz9H5qB5eZCPmJDeO9x6tgDdEA9Li+HpwAtgpDN5m7BNQ7/JKsP711ddPJmlqdS2vQ/9GeVVQSFi
WxD9+81qJzZcOC04GgskhDkA/LhJ0i0fkc+XfW3LwAdtMsPg1/OmKFA9hvCHYf58L6gBt3uUpQPW
z7iQ/3irnl+dZ+VfBUFg2vBqsVfk6chWhuLV2eEcozsoKFByDMFpMYgFLJ/rGU+6C+Xgubi6Jsq+
TvvoR8yPzw3K5S69KNesxnOyM67ZUBImB01k33AIVS27AE3M7uGkPUuCo1N8142js9uyVzPC2w4c
7JdE7O1MKDbSRy844BVWrTPhfkPKXPqKOjKMtIhX+ZQxF9gfPmFKvzvKFH7qvbk6ijxwif7qo3lH
0U8ym4LXagtyOoyjQ0aQ8ef31vfUBIt88pUys+Ufo4UP2MZWOLlTh7GBeq3/8ONxKTgFHhoKQWcc
nV5LWWh9/HrN793uZ55Oil+7dedgYIYVcV8VQy5d0ATZZTAAczjFxFFA91P/FZjTm3Q0wpYKRy8u
jeWZQ6a0YePDaE1b3dcUGNq2BeHg1Qbofc/s+im/0T4pHWq6/sgZqnVMg6aQ4EQdFOLT6ZFCatDn
rIxdO/k0cGsFGh4F1E2snwr8NJCt5OZ+jFio2Ij6HMAEXJrjX4NHL+NlfE9llbOJEbwcFrvSHV0C
pkgyGKowMU6NSrM6bE1RApDZrFUk54w28TReAbIv9xITUHBrbokjlPcxnRBJ+9HDrn8FBtK339dV
iR7ri/iffO1TWs4OXDXPpYV1xjzK7j1Q5z6tX1DZ5bUXRHa4oqGQ1uukzPE1zVwiHOW18z8ZqySs
sgpAaWNdm6/1gGS5s3fsz9qzpVAqpAONQwV07hC+WUt7CkxZEYuEZiYMLZY6o1bjMGGId5TrGQlv
Nkde5MXN3ONKEnrheuieRHd0FJ9NR4lxVQoRAMCzLNItarqogbj2I3BrP0Yd97wksd03KrGbGj4n
GTgttbGzvuKt/LxEtt/w4dv+gTTMP0Ybn4/8ZbAW7AEFmjo2chDR9W629uiucBHv1C5JAnUDY9Bb
GAjhOuYE7DadtrU4PYlKVYZb5tN0TGdotqM6hOFeOAjfBJgwpHvkumM2XlsP5o74wkXiosaTr9LT
aztl0JuajOeeCILWpHEq9OPKAmsNuz9yz8CzOi19HpH1hS9h8sL+23XDxL0/F9AyhkrUpEfC6Cnp
yn9EnqhXsL6QnjaMGu34fUn255EwnX4in83ggaVRWyvy2ek38tNZdj0tjAuwDcY0ueTyGNVXE/9E
J7FUOTlS4KrmDVYJ8M+/YgXg8dwfL64vM7UJsJfak2ZziOGUyqqoct08op8J7X/GFqyysqnFiHV1
DoPe64Mnyu5ZByRsv+MJe5ihtg8eBecTqx+FRbbEmSEcm56BI0FCgkGvcflOzOS9QW3fVMlypMo1
yU/C4tQp4fynLpfWZqgcZed/KgVwQ+hFXHZOVKyquEkGnpe6dE7ZJzBgzX8o2ZyccEHS3K4RuF0Y
H31HVvWXt91ad24zmSJz1PwHYpuAAw47fd35540cokhHzFloB9SrF2sMPflHK7l5HrwZb66VRcHV
exb37ynmo8jZYkma/eWBIC9Q+0KYa3rYBmNHd4Nd9/+/ZvoG/2hftOOpFxr001o5jh4/YQHMrRax
vzJrzAtdmm9lROivh5lOkVec3sMTsX+NCdYg+sXLeCHTu5Xj3gsJ5eVDx5wljZ8ZAAdEXdP89ROX
0M/hXeOPq5LXBGPlZi3yO8Nz5xs861TLjMCa60YlNzL/OrfFSaWjzSOgASXrw1qFjycXo+iE3+oa
p3GQ0kU5OSEol6lrh/GTTD/bV29iDuTBUccUaORm03vw5bgMdwgpXIEOOUvaMcsMW5PbwXsVUcO+
yhhuRVtE1oZF3Gu4lSYod8o9N+bKMTcTPgQYlbntuyEYjLqbjWAHdEz1/PjzGMqu5Xbgk5zIuxjt
qkaH6YxqZ/KKsdisQblYfWnsg6f4yYat90ak5obJu5Kp9kbihw2sj2Z1tbPZ3xWKWamLQ5Nr2c2Z
i5nRIfepW88+fJhpMmSXiwb6OKtXO5hU6CzKknOwW1Zu7nUqqjGYuedC4wcjVQymhph1hRzbyhUQ
5ADnQW2IgUdyWo6BhnRAYNUA8qoaqa8s1pw860l1OyTXEKoVTkZdNKb74abwllYPIBotVaY7nadP
j61y3R/UXGsgoPShhSy5DT/K3UnTQN0O99fiHMlj/KygqWbSSC8FEDWAahwBUYCeK8lPfrSknrKL
KZNDZoTscm9nZ5VhSi2k77i1JgsEgVFyV9/ntv5T7FpHqMvHotmvw5AEx/g2qml1kzm6/W0FlGL7
zQUyeoAhIziBN9KKUvJAegA+IfxkYyTQCJBBkdfnQmc0KmkHQFPgDRBUcGfexLM33hL4qr/T0rMv
qtd+9jzsU57SjHfFab3kxUStNH22bnrhIsAVe9TQVklHBqhRRBclFpksvbqKqD/4R3Wt+tdw3HvN
zf7TnATOSxkcvI4MDdL2YYTKCtiesTDbzdFJYfx8wKgKD3RQ3HYi1w4dMlLQX8kt/s+ajAIuYdC4
Pz2657Mek5UhG7pzjA9R7MaselmBOdlZTjEZYIBnLQJH1rkx5EFl88xbb9Repz1zfS1hzJF3OXl0
LKidzewEn7pClYB1kN2oX+IO2iC8LuHEDgUfJdo4j3SbF9pd8h7P+geC3B5hwU/r8h6axQIgGdEx
M5Jll2/hUS9h1xkJl7xDrKn6BfIuhdpVVMvIqbxKw460V4JkTK/55TXXlWExgeL3X2mLQmy0+J6e
7xd5ETi6ls0V+z3BarkgRXETctul9miBUdJA7cLhVYvlLY+1rCpNO2jNZp2AWer3fB1NjLGiTykV
cgTUlUbAbYXAHdJfOxqoUZfnq7/OeFcp4DMkJsSCJoeYTUJeUO6gC1azx1CYz+Kj/JL/JgMCEeLN
gRbzyJoeFUr0pYrfZV/0MwLTxYdWN/+umLWCv3Meox+e7sl1WmIq4dJvAFDOWizKgPCY80LQYZOk
tu4ae3DuzaXEnwDILPCWDvBK41YSpx8n6iO07LaWMBnLKDMNVMfAMB0UV102xpjj+w66jEMmq7fq
fLQdDazVALxDuCJ5BbKETsOivrL947NPUFSHfG73YirNEHqH3GLTzuMovSh0+EiEqwYHs5C+xbJn
1GVjB4ut7JmYY5zLCOUzPvI6O4U9/i6/66TUe+Vf9aqHk6z7Fb9Gv43Z9UrIEo96chNLC7207j77
da4lmmnKerni6OpnTBsr1MekEq1TmSxiirxqRgpRvKvDNiC8gfsjQCmb0AoCZ3SL/h/roUsj8uxO
r+7043BKBvPRa6qN14gE1LgFW/ZPXiO40Zfnk8dHWkPsPALO5Ukymb7YcjS0682gt2dHSgNG622M
V0C1a/0gcno8HNP6pcA7fSMO1qP8y4qPmXBIaRCqFH/pNlP19AUtIYnVI9TPJSc4DsLkVLgb4x4t
T0mu24Cs5+kFa2lVyOxAT/C9qOvTwDWjZ3Xq2DjzApwVzUc716/tH2tgAhAIgPek7Yg4RnXdeSEC
Z2a+xWM81mtCfF/Vphsv1KHgpb4xbJEY33YaopEwSkJu5Zjx1sJZzo12CDZhyAD/w916ISzZM0kz
vqM3O6F5aNlY0LCYsbgxeSFf49EgwREk6gOiiOcFgj0+acDgZpt+mu6Oc7YKLNUAUxMnkKCxyOJY
DwVuwW2U7Y+DP/EMg7pK3FC7sUD7gqFcRqSAkzxJDy/UZ+4t+B33tPHXxwQe+g1b6YGR1OmPd4Xa
ImRoK1n7xiJsbU/cV8k4mkYz8ffUXfUrQqmeaKel84EBOQQauoFzxITGmuXEaH3tmCsRKFVEXEni
+mCQHWuPlexr0Yl0+Z5L+QtDu1XGbR3v0lU1ZfVyTsjeAmApf8JFNh06jYTTjLPS9MPyA4MMLu6W
sRCNxLw5eDi/tvIbSCGHAzSBdv4xkkFuRuz7KaEuDG/mtvhi2VsOAGDg7ja6WXzlTucE4XMR2JpG
R7rSTPmJ8KdjgwpXSMf8BB0m6vDj4Loygic5Ua5CJ5+gEJ9I9eoAv8Kl9BjoJE4zfsQzDewYHeSt
69/nwn3gOvNkfV1A1ViIw5VV71XeZyn/YXwcwx27DkByLPGbbIZrWLM2yLuEMLl7RSkgQ8grYjro
ZZjxUQlIiWDHxiolCkVaK4eJHK1FG1V6EpE+XAL9KBoN0NfVNTeNbAVHaM/pBB05jCph8+4TLfu9
yJrR+/CUmE3LAfCer6JnkKdZiqGXw11a3uBtp8HZD1w+sNj3d4Eh7Fg3vtRIxYingjQZzK+liC5S
BXaihM73fqRc3Xe61LcXj3sOiNs6IwWDHDMG+OlOj5hGs0mWHXQGoQizfbjOYFjbQrPkmZZ7Y37a
88t7nYZIbk4CkyhQVqQf4zMcGR0hxwfmh1A5GXhDZlV0sLG0GeaVNbNhNOdtQmYalPu5gpp7rkhY
mizoWU3yQ8SaToOEZ831oIhO6T2czhTzLFVsZEdkCY2R0PT2Tz7AWL45iFWrT5mVuuyCpgQq0PXP
tHpXqVCLMMeqV90civD6Byp+6YwHowsW0E5jTKp0KNNI6uTw36aGRtZEyMsBEjSt6+qBWqQ6w8v+
lz1Gy9d54n43/Ab0CtVyyRft6rG4c9N84T5eJHG/NZ0OQQ4vUIkW/CKefI7jzR6E00nrq/gIEuaN
Qx9qkGqTgaFToEVmcTX1hcXz0NlD4fb74iaFP3FjpWh6bwGo4JgJk8+pAASAWH4wC24vAUUtI6gx
pXhrvbxi/OI0GI0J0OWHuniuCLRhQmgu2I3y2nEpp6PemgHAYi51hOYdhzTPEMuTs/NrvnpH+Bou
GbI4U9zjVABFkcu0/DNqDitKb0EVur56CffRqeaZMpRapy7eFb1HUDh8B8QVsf7ZfzrXnEhoUIO1
ZhPrq4DbIO8Ed3HW1DXlDCKc9S4UlMUl5yjH18AYWk5O58hfZJ7tSR2BX7kWcNzOnus2VMifLkU7
GwqMxCBTaPsj6iKEdlMEylP6Pxbh1mirmm2Jjcr3SXK7uEp/Oe3u48C4Rl2LzK/r8RYvS6STeggE
KoBZYFgAD91W+a774njYIZy1eDmp5/5GdNsYtgf4VS/6XCS5//aXaIn7IuZxZwnq5Oss7OuBVKGO
+uXzvn3FtYby7ZxFYDCIFHbyu1wYnOpKmQz2/8uAGZoeq9vei61IVM7WtnAFGusQ0ZpXjX38wNu5
OG30Ngp81xHCkiLYYL6UKbJ1ajvoxE/uuDHL7GQ5d0ZAIoyJDLA07xkKpIdBXtzgZAyRjbRkrVYc
B+hsSDWUa9VvMCHRI23dQNt9MchaSKSJmIknQnHWY8hGyR5ufWvBnuKIHO9xROACOR9Vw3Tvp8cK
Gr7MtyR+TGaXfwcJZBl20SAhj4AiQFKX2Qhdu2f9J3tJ6wn/lvNvFbUAmJWoLuFzHPMl3zYiiZfp
zC0i/ehkaY16Obv5gfs1AuDc1NLH4PgrucE64WcYgaIWCxdEntyB9ycWzEFFzuKVgue0jaISAnKq
8iafwyqLNLbHFXobK9dfqFzSmoFS7kTSmIwc4Rlmau2kUlvdjJ1fn/4UFSu6fVXL72OqK4B17bo3
nBuVrRpovX94tR0J/tI2xe7BjCCDx76SVOrtAVcLpGt/ujI14pEslmQ5spLFgOs1lBK9ctIyM1tP
5w2eizfu587BOPZ/467YQCdhNFznEDhLDBj2yCQyObRpTY4SH8fqTEX9muG2gucbN+m55HawkFEM
cGKylcKxlLgRI8VOWqxGP2WXw0TDBGwyBW2DZdjeLWFXzkeuFaXsYUcsrOUZ1eslGgOtGZ+0wC4E
BeTbMQQBSyW2y56uAauJuvYBFmVs7qvYD5wjaEKXUqJBbT808G1pfAO609QHefKdouxN0PWd1+sO
czL4a5tQIYc+a/LrbOsBALfRniR0MRpdWIQqTR43TdyUgRXW9rkahi2KQE5/3ndAPBJBniJWJKYa
GDOf9OrcoBYKnzmSYPm2MAUTkjZup+ZIk+AiUWtgRHCtRbaXRjXzIEU1FVmkpUJBq8GyTk+PWv6v
BIRAj6XFEr34X5Qn9WPW+gadRehiFfcJ1VkPzxCZdnJLa9oyIAsipKOavOiqgC3kYbjCp7GESoMo
22zpUq97f7AxuYD/CSO79hX9SpOkd5cVy753Z7QE0amO7EzNhLapub4xxfUxbkFWN4lAwleERShl
TnX1hhfB0oDRykdkAy0a+xqbJzuJCXdhWhLjlYK8f8aZXEX9uVXsJ/iZcMq3GZ/LnTwOcw/VIurF
hie1mkYZjrH++/4nhpMJQG1kIUTjGYeEgnqVhwKkyHe41iqMq6XLSyYqmNavUD+gu39WBpZ2gQ/U
dpK4YXUVBQsfFvywOplyYo1Sq1bD/N3ClUJ0g8JXtyyqbqG56bmVD5kn8U6XQDaw1cvVBpqpwhNc
9HcRn9zSXr4iZEq5s+Yf3CjtLruSrNKE0bMM9nPbIgURyTeUyqkj91XK0szafC0oAM6ZUFyQoqrb
o15jEbvSICpOMgRkpRbzgPIzbeC/e5sKX1MTldRi+Z3dLAONZmAEYGO3Wv6ZDk+jGWlSOFE8yR1+
3HEW6XQe01uf/+ElMp/yAo7fObSgjPJdbFTcQ0evnyAbZ05wsjo6Pq1UvZL9eY7aVIZD03OkkQox
yBAukZ9KZSjwv6MP2X+USw8Mi5hrZCI8eHrrtIpwpURhDMYqnCkWMrvUKjB9APXQva//pEWAy5RO
MlLDbmgOz+jWpgAGT4EFCgp395EUEoY5hyMnv7H3KOo9Gr8cbp8E+7NQj8VlG2GKlynSFFXZTfr/
m1PhsUXPAVHELh98Lx4r7BocFsLpPIlDO39mnOaA1a5X3MoQ4fm6Sf4o/UNOCmMi9YJ2XwfiopYo
SP/z9s3jLKasu3SJB+GIAD7am/KapncrBjZntZKr53pbyMgXpDihc3UG1TMbsIv6ppBDTUoPoIEu
Qn9n55GbINDsG+ahBVt04gpZzKQx0NTFmfPyRQfIEdMKojiZceOSbd8ojFw9IMu4mjfgRQgD197H
UVWa/+p4tm4ArUZnNThWicnUhyNdbV3h+A82qU803Hvxwc/ZhphIOyLKxdvpWylxaJPpmn1S0qav
WHIF7bfv9iWbnuPPoVORLolBetV/Zn6pXsqvKAAQ6OfhBILBGJ3HyqPJq4k0azyNbfIFMD7eH73p
zOocE29LRklZvBGUfQKFmbu8CFXcWemaakeKpxvVJx+IHjXKoTZJ2cQtGyzsqMXqhn4oscFtqdMH
eyL+KMH5mZi11d/6tpXkLlUBmXWytI3Eisy6C7wGZgGWutS1VaM864FG4byLRIgI2d2f2p9KW6PR
PvavoqmpqWONEvk9qa4R19SazMbRKWpBfgxkjEXwaI7ZJ+8zVzUnYiK5Lk2razBibB3JDy5AxnHQ
AOp6iNzsdNOTGNjZjagYjkwF6pNWWbKa2uUhyxhn4SynVYy4rsV8cald455CkHDiseuLhcsEXNwY
Jb5pmYK3ca4fhBxR6JXdVH+j+fauAicvgqfiai0CvGW2t1+oYD8kQCaWdugnI7Bs5BvUvPZ4s0sv
8rZXulci8VHzXttXwZRLlXArXJaeWQsZWXWFC7HDOJuqdmsaXBVJMfZueW4BvGSYH21dgEpnXYVN
/I9qnxWqQk1Hj/fwZMCl1qCrZn1N9urneHFdInlU3gb9vf6EiTc949gviP5M3LgTeViWiqYHq9YK
NmhJ6wysxR/S+wkLew9/UNW3xi9/MEeVbsHdObfTu+r5gP8nFu8/LFoeGZHWL/0Dk8jSwJtvgzej
jS5a8LwoHcCBnD8kLaM/Psb6ecBrAv5v3AhQELKiw9Wgm8Bwk28EE22qgx6FslQXOj5dCQn90hoy
+BQFp+NGsjj/hzRZXR8kFFr/8KxmCDc6YOFmCXMKVxo2HY4K+CGwqjXZz2OEuhp4JKnXLMJRQV5w
AA2sNKsgc2H+0j8zFh4Zuo/jZMxCdidp1GXoseHBzrnSLaORcQBtCKZKkMSsrZSlKNqHlnGnOuX6
/yltq9Jbqo9PYoW+6gGjQ79mE4WiIlZ7SHdBMmGdyfJTqQEJ7oTSgLmBKrNpDKNlUFguSx10J4iv
uHNE4NtFg+0mNeGE07biA/EqLBqpVKVtP+2ttT5QR6/KebmichBW2/sqZj18KKu3xtJ4kzqhxrXI
toKpIDwYP7TqbVHbpy1HfAwxbIH1kOpyChOIHk8XLvLStK+Ql9zvyUsoVYA9d2xcr0zGWs5LxFYK
DLH0PdA1Byj4oHKshAOGO0STgfdv02uiRRJ11leuAg6HQGzzEdUS6L6E4NeR1RdvXfHu7HEanucE
ZxspCnxpJsaAcqGcZUVJr8I0gIyFHU1XVjlRaFw3b+etOEte/GpTMucezxRCQUOUA5BiRw1CCgoi
fotPvHLSfqiAtNdaCuzkLkd+PhRnuXYABIFOgSeDwJbOpw+ki+6L5++ck3znafnq5IHMqYnB9gBh
81Cy/zaDCJ7JnpNa9CXhdzOJpwy4LXS/6RAepXyTD8/HXppzSRT9FllSnBbkkihQoQ4YM4SwtnAU
/K6DJsRUMzm2kKd4fGRUoeMwLRvcvxCcGvQIyPyckHrm0Nv2oIvSKyysSOdGPF7iy36NXJHVsp81
wwm0uvgMENWi9CKDqmJU/nGGkjr1OWQ0VBISdIrIsJaM4RxWpUGs2VZITxyu+Bp56mq65QjYRDXD
w8SVrGU4dhmOARahrXgTAZxptAnyFzHnmiwR8lsyl+x1qMLVUHGUPtrP3Lat7biofx7MVbqcAddU
4DzON/K5zoLGWQywwVJnrD7e1/Zeh4JsEo92ZMMJdDz0yAxzkYj/dBY/DILWc6QkhUayP+kkJsID
zOfSdv/i+BqqKtciylEuCzcLJJ7lYlaPQ/w7UGTYy94A50j/bdQuXJ+vBDAKxTe1/6yFN+Gxl5/p
Co2DGMuTlYQ0bUwKPlKI3TZlrWLXvHGi0PWXlMaNDuIV/iMJ+vWJm9hQP5g3323FKAp5e/GJg49o
FVrVnqm2hjWvW7Mpfw/t7yWEBdpPM8FD4SdmfMssrB2dO4ESzoJxwCpVjUESfF1RyWrjtep/hf8W
Lro3YGU+FK0Fk2FIWunPRG3tx+1tu8PnJjgt8WxWoJsEfi31nyb7mb/yId4PzKC1iZfZwqAzyjFS
KhgIM0YN7J4p0FjzV9YUEm/NqGF82Hdkcs0PzMxumstTah+fBc7E1fbaFyLee84huMmGCmrhj1x5
7kq0nBxF6skVNLyuteHjY+l/q30bkYEasHzSPfzKjv0uIiNBGfPSWFIpVz85GGRCUoQA+TQs7Tdl
RsrNQ4ZuHLVvyqoFQp6m8xL6uaYJdBpWlRnzeIBGbn+v1S3DxKeQOZWjVp+JS9Casfjkl8rcyw/L
R4RyVz/k3Hvof0mjo06jRb5jj3maUjAtehxy6qjheS0W+eq4ow5D4KfkOOmWvuajXx1YhKR5teEt
jaYDDqh0UoNVwo5FFT6YrKiT4gw8c97r9ZIHQTwyZIIYbszUXxFpHnoV6S/IDn9KobvpYJM6ldJT
KB9lvhDeOGoc7UuQ2ZKHPFoE+iEjYROkWYvp2F9ZRlfGSAeIN8Hoii6ym5BDLvGkgsX5MlTLwBPb
oP+QR32cajxCn2xKyyeO1awiDLq1KVfr1v9in21LK6otSXZSHQQTJeD0RkQ6WXZfQafIH2tmhS34
NWIgfg2+M3CpvQAjnR7YGPThBUs/UsmNfASMdQ8whuaL3yIENa3Z01PoyImfBoc4Nd/724+wTy5E
EpkOTIMOERAEbtiP0zKUly29HL15VfqForCf/hiiO2Dtu1QIS5+jnl5CKtgIgTTt1oMMJt22p79G
Rlro3eRs7OhtAR6NKxVnAj3n+hNAMw8/x3qkC4zCu8SFa6Lzgxn2zfadiaiJCCx59pPj8UqmTte7
vAPn4eqSv4kwud+O5XYlWScqSXi/C1894T7eV+vpPDmzuCpxWnNKOX86DGlrqaI6PrJgCGSndTvk
RubITgrIvn6T/xyPhJpAmtFWlIbF8dJfQmKpYnMMLRBNvTxL67FAs9DWnAKE38VIoKKx9gZyvkbM
swAvKZ4LDy4OEtT4BX/7g6W4Y7fhedFozPeNJ8Tx/uDJdQRVz1r0dGhZ4yoouXT1neTt8DlTWHTX
IP/kWuuMNLfeigIfdzVJPqZSxq0XvDU3R499R1J1/rC613TkS1UXoDgnjFXdxyPxroWonbod7JxP
qdAMlI2l1vauvfLIQsDbKES55NSsdCVPHzI3I6lA9UCAAPYl8q05MKzKGtDAYrJ7yrDs1+74+P4j
K7T4zd6hIoUWwkdmXAre8fr/+xVhBuVNZ+gXvECUmmBcpuIFz2cWBxXCI7vYhB5mh4WaKGJF5QV5
EzALqHVFkSnTdWVa1/k/GhXlOa7vlDF2Gj1c0JlwKnsg1lrNLSJnVvKGSx4xYfMPPiLXqeb8IcxK
6PWLOclHCvjI8JG6pw94zFeLGyTVYpRSfCGSlOFtzLdIskU36OlpgSAgoC3lj6cZ4gg3uMqIG4Sb
RfmJO9lhzapaCOtMjc9wBr+wcsjzAaimtKkX9epeo4jtESzRrmNPLYyDJ4vDur6lZtnymc66axdY
DdIE2KBpumVVgzTfdqw8eYRU8Acqbz+goHNLxr0wkWbVje4bvmLrzjGuz5D/ciwhTeak3yB4IZLK
++dby84dRLS1eIs6EliFwTMkR0oJ9nfa1hooxYV8rJB1W8PfnJXngOr4opXIcCjgC6LmVuav90cD
YWrEhAxJBS8/4dmSb+hxajD90gZjBcE46bksCk+gX1AXCLbkW+r/YTC2qEDQtAWDFKCfTZfBAze4
yMlHbjMh8N4hp96W0xrhi7j8N2qMTgMqQVfOCr1rLPZJqVO/6Nf2C8Igy5mZN4Rj5IdhKCrPqblT
6en1VioA/+26yCr3rZpldpJQvRi0R2Fk0RBuFui3uX/jnVnmLAOAx6Rkd8Blot3o8r2t4ngEDl2D
8g4rLPXm3duaWdbNgbx+hJD8YliXoUZpfQh0PmCVrlDDs/NpJ2at1LjC7TaxWPwYS7ojAvAJLpGl
OvOOYyOQilieXCWZqusd/eL5q7ag8XCZDRdZt3qopEsgvMLFAAQtplF8nbJX1BYufT+jCSYowYSO
pmoHp9mpE0TjBtmn+EQZ5fe0ptDSMT4mERqMsLXR3yQAt0bijYmanJUfwSD9lGfFJ4ijPVjl+g4l
IcTAxaiyMU32b3AL4D61yQDiX9KXEyLRhNSr4lXXBXlscu+fNn8SmPUbRylIzF2JBRIFB+7NAuks
OvAYAE61C12cCEiue3RBm3FyKyVYHn0d80huzXgxfrLUpfhzw5aRMB6u1+OUv2l/6NMfsJfBpHiN
MFo/OxR0SVqabxg28YcsAuhWwAvsBj6oRLilqsOyjjIcr+L6iwUCPSb/DIhVnhCWWQLBnfvNXfGM
o/dj74lF1bKYGqZo+mJ0pxoPJwmkf3MHu0fDI+PE0W61M+v3/2/OFBM3jtdFzlNof6WFpKsctIjW
MPPGuFg0OceEmbSL8LoYuWMbOwswq563DduYV0ogmsCLrIDyuJ+stvhoWuriwIz0SJpiGSM4WAnX
w02MG7KeAqMk75M95T6LJyDK6dd/2YIav+17Y4/XwZLAGFFskis7FBEP1oEgm/TRwi9zTkqm4Llt
MNxgfGKaZhI7q9uoOGYjKULpDng6KSiWwi1FiA4Jm1eqB8YhkM18AZcGK2gwrIyLRaVn9bRuuNTj
i0+/z9sJGFGev9OXelfXLAFIqUHX/dcu9jb49p2PZkuDalZOPohRdwiXpCYg1zD4UmnBz7ymqbbQ
rB4AlwSENHh4EiepbOYBKLcy5n4An3o8D/GqBY1BSGyHmFOjmKnqGn/tF1w++foiBTfYiSoHC45j
iFhbO78Q5EA/Dce8A7glcQliZXNxMeQVvb5D01fB/UZsyRmbHwQkHqUpY9macgiyXXOLh2wbjZHP
VEInqkZYLw3f4coBasa1JzLhUl6JmOb2WUa0RKYvh6L1CHGpp4hGNOoU1aWu5aX4nrNqgQdt6Uiv
E7bZvC7lGuUE2/C3GZ2cz4iME2Gh95Fjjs6CE7W35A9jVqMQ1UCRPzXlscSXOWiYW4KNn+wsL7gT
OBdP1T1N/QH8tPHb+7FEdT6L6vA24rjTNiU4Na5GFE0Hw/uol2r8pJybBM83lZZFGBKnkQHY+MGR
uyeCzMnqlPxFmhgbO7WQoyZg1y+zrFxutBvB9XeNyK9ZwrPPs8m6OBrNjlIweqqGXOU1mmh4uRCu
5G+4iEnV3crSuuJwJCSpB8zOAJsu3Rz/6wonZOBJMpxV4IOCHJb9eMBIiYfNq2//aadnlLBkgbHG
/VaWpqmk8kp5xnHgZj22QuLjVI/iZQLE7LLSEQWxkhAge9U9q3/+jVC4ii8YtdQCPdNj64eFqhJ1
pp3tDtuxE0ygOPL6UyqXv6L7CC6KBlx7UWpuOH7FOrCvbu2hXQCPkK9GgMm2pHKfCbeAojK+UvdF
C605x6t+am5w/HOGrbD9veD/ktRUiluv2tC8/i5hqhwXJ0dqtQ21G63EVa3j4Exzb06Zr5rb8tSx
IqKU4gfsAlsqwjEofK7Gw3h44HsISu0OHAo260JJhQIgzVvgG9mE09anv7/qvsVLGjInDLvl9869
+5HTmEJlq9SSU6WrJJrko/oNsp1uVJk+VUiMEIb85RTI4PgtisG/8Gm8RMjtj+mPRmP5mF5SN2kP
BTfeDcr/YlCTRkc/BpCcTEkId/n9VLzjfpUpR1O0d2x/qO3eM1DqNUm6pzs7BM1kyYfLJmSjsW9+
+O41wgJjdn+xSChs38+ng1ZocrwrazacwlwKjVRARBu5B+QtrBBVQPMW21gaehUmK6nXabb060P7
g2dk191sFZlRAWV0o5kPlDMe5Gm0M1a/AHP58HsIjegIggWMUkQ5PI/jfSpwQK4cOsKyrSjngsii
XrLBk7yUrHwFhINCjC4okdRwkU3cVqLfzMY/vzRmXZoQwu0VxRStqFiNabY+2qvgeojC+ZJtDkCX
VuYMIlRQvyy0DtRTc/CheyVZfJRecaR04dKELCoVqpLPiP54aJjBgXdAccYR8oFyTZ4Rp+O8oelc
/1GnkHGyJJBqA4lUNKM75Kd76h/lNtIe4/07I5KyQ4UIoKaaURjGppodLYpuwVujWWonUzuW+Su/
0ID7mSdZ3j0+7TqzzbApJ219W+HAfldXrtDaWc39uNiP1yraLfiiyclzBkqav/Hb+XVSuwaZBsJc
2838pbzbsqM0Tr8ZNTHYtZ1U5Yw7ZcNaA5JKfAJY/WRBQT8y4PXxG3WavAj+UhF7eHFgpM4ApCIz
lPaxXGCfO7e640rYw8xNqL4n/+2syh0wk93BfHjYLCqf/D2wRVRPwc16DMoWb7PeEHp1T+bhkfjL
c7gOCA+1qjJU1D+M6wLL7FAPpLSpFk6LZ7s40sEQJMSgCfXEHwulcTSqNPGpHGMcSPg0CYOA2BWC
u/uyP+snxtolGMkETX3cuf3dkAqB6SDDwJI/BlWRC49kB++pfQm/Dyp1suWDklWK3YyzlrZTA89j
yoUlYhPzuuMcLOvEQ15gn2T9iiKFwaGoMJGYFe1Ikg5FFSbUMEJgl/j3bQfndmm3XMDs1L9bqHMW
O1nVuV25u7Atu/aE3pEfyHPKjdprOZvbfydXWALSptHmTDz5TN0dgX7dRlMwWYGyrN/AjD9Pg//V
hN9G9mkiLODuTJvJNXif4Mu17xXCybx+7yiM/AsMTZhcJtcTMsgKG1tv9XolS8soG8wHzJcX3jMb
zoblmGEoI9RCv4RYHup9RJJSSeaPnaP+lHoCOAZkXYVIBdVG9jRMYeTsuRux1baDBXOKlLE+nb4H
6g3pAscsl/Y9Q14rhhFW1gRvBIE1K2etAF+QD5yqJVsvltlnesxT7qkQQdMxvCIwAT4I695Pu4E6
rKMs6/SNxG8pRZGlcdntROnRXoJL8kS9EXbYFgrBrGiRNhSGjqjAVOGT8rPMQcdIpV3DFpx+xDGf
JmjQA81qOsYVBdPfbZEMaUz5oR9PI2gMrnhKsrkZN0V9XM+N5xdyak/Dkq7F9cUo6+fWTVQIWO41
6k5A5BIssIOF60rh/YBbI6k2MERkgXfwO64S64+KeNsIcDcChlosxssQNb28XahUJpXTzyi9BaYJ
hxkVHgKnbLIbgIaxmkVY4oGhSTI7UiMkc5jwlupU2ZcMXjx9cl9dm2xyAnPo1OzhUXxPAhbyQpY7
BedZeu3Pjgceyajd3ojGka8QCnSxxeDJx769pQHvOmJyd5HWKocl8koq6XwbozNRAZ8gFEEKA7a7
+5F3+6TmYJlwM+6z3BpCH0C/pGL/KDqc/bCzI3kAz86noH2mmpJpdlfy40rdNthvBlrFMUqCRmXd
rkbQGmHmM4zGqVbHqIjm0vX9i8YUHoKcsSq0yyd+YMD9PoiFDGMxL64Z31PannPW//yTKueq3rA6
3oH0J7eZUOSMbkqvkQGS8TF61ByIkL181Uy2LIA7mhbvSS4EC8PJYkmIrRorFV6eeCzHTrcTIuvu
Ve0tfe2woNG6HUHtKc/aQn+3/DkrkimIThHMTViQ0Jstn8W/ueuiRdXOs9TptJoMhq9uxPqeA9tG
z52AjpdyZ0cvaV1xq8HY7JPGC0+nJ5JBsjV0uSipTQUgTNIuVpbpIgSb9uk4JETiEyFOAlIbQ1AQ
PsLrQR/gdx+7QIjVMmvcu5Vg3yg847r30W3nn5rlI1PitjGdWXldPWt8pE+SYHYJ/eyuwodl8YEW
OkD44YDWGiRGPSuF8X7ztG8kQ7CmNSZvRIqSnzhJSvLrMB4bMIzoZoBzijFamxV+covRbyDdV1dh
iz3F/NLVSwPLIz8qT4Et6ZohPGW/06LNdShjvkz/0F7NI0Frr06vMxAb3p4o1lwyYluXSRqu6qMJ
mlTy/XH9B0zFJtQUdJUPy0DiCciKJbJVIjwlfiOys2+2h5oca8xRRPY4T97PRUMGvwg9ok11Avx/
gvQvtZ8bcsdzqY0ZrqGK3zQ9Alu3MiqrYmT+sEOpgFFIUgGKeCyn4Mz+Hnu2kT70WbM7/M3+fs1X
5MLHsaBNaTIkBi9i1z2TZke2nZeDTl18YMcjaEpIhAIPUylLDs6yOaNiEZQoSQnKvx8UA8ZZetjl
s1idyvpTbp8TaeUmr4ScSwYS1rBhO/XxE50FZ0BJJg3iSp+jV1zGtaLRmHJUz1vs9KeJSycUtl4B
k0lX4aTZVOsSQJOB2fHUEoiAMdUnCrLfN+UU1DwB/VLyGObuiJxflAhtY7K3ti4HnuX/rc0y4HP0
0thlcQ0O/hDeSzdi/LZLSS3lM+V2w2I/XGI9PK10FF4OeEdPRhLuYoUNuWfUO+XOsniVr00u5FYB
gGmb1MwkH8O9yGgK87x5LbQSqA8OcBwlAmFJ9krOsbO1x6IdmTYeGKUqJp22w8AjUqP+PsFg/M/k
h8/QCkjBYH0Q4ip4rSW//9+MPmOQNwaVcX6u3wEjYKSteKh1d0MrMcs22zGCJIVDe9UIgN9rPb4u
G9r9cPG8oxX0UYiA1i6/3+QJxLhbTSEYYfjst9Og/NgOi7S7V6oAx5bauzTuA4XpkKYq80kBymTy
sCJu6gcqk+N0MtK8PphanUQirnd0y3RnlHpDFeBRkm8SVRcQOsrQofh2jGPXrB3Hh2OATuomIHcp
o2q1NvpMDWUORn1cN+UJ85C9bWQC98fGfln+Xgzt+s/Lbj9cyByVP0tdpCbyJ17+WSBZPFO8Yh38
ZF8GN8DG56YG7inD2E0O7lRbGFfbSDYapSKub4rp7nL5PAXRg3CtLTsPFuZpFCOj6uuWq6x2T3mL
e33ec2Un+Q0lMp+1ckVGjHh2MKvG5ly9yG3yCuQ1ZSrI+npBJAZEpV6UG7OFdLz8JqBwO9QutTQm
jzRY31BC+LKJ/UFdCoj5bi9JUbw1m54X7LCcPg82NZvmepqRE6btVVBWUrq5wSKAkjoCXVW/V49O
t5tq/NWggP+yygAlK7+Mzz+KulmtplMjVsnt0NONegOqh3mdmPhFlZ+cLZ1Z+8i7RRs3wNI6Ik1M
uLVbkqp1AoCnt0ipa4wBE9SG7HMCXz6OQZOBrMsXzIpaRYl9Zl5pvtPGK78ovvJGNBLK6aWqeFAJ
AlH1auj964hVFJ/xW5UkfrYZwO/DKnQ8+A10zmVObVqnhqR0K8au1E2JHXIeIxHyo2qCZrF+8Bjv
3lDHU1l1KcxZjMC991Kce+6rKFPwbDp49oGKRqk6nXeIkjfEnlwzn42mZVbC0GjfyOpbTVmFSWnC
QLI32Wy0LQyMlf41lSaRKPmTTCicWaHY5LDY96TRcUwxw2ziSu3CIRU0SsbClMQMp3NL7ki7lvFz
3+NyNb/S55aVAUJWDG6AVhGnWxP4joXOvB4RLVhIBFF9p40BC1iMWxfkI1XOAXFNh6k5ZiKSkZ6T
oea4mrKhenoP8PtGx5HB2k+IH0RoTAkBxum4MDtigjJ6Ef6dacwuFRLtFEoE1TrcNxXh7jfr/n6/
vRbpxg22PsDNvjfyr5Ufb+iu0nB+ZOe+cxa+Oa5+JlTTUpze91fMSM5AFefDmGKyV9YwXALPVnSh
pG0gV6vZ+OZvTbvSEnq5ZnDuOxzsCNUOSMBZ3vA9dSAU+4wjaOE9carPhaCLPQbBp7tOicEEggZ6
p38aOzotmK/ClQQOZ+wMKrmoZrd+CgiUxfRS6m4Bp6VLcUG9qMRAKA/8LpQo7Wo5MJZycaiVdclI
sIvt1oSnXyHvKjA+i9LeBU+Mfp8LTtIQWf9rbNQ9vt9GEZfQwSBY3XaTcW+PFbp+oZI+VKaiOyKA
Q05d011Rwji/sPpImuWRvy6uQ9MUfs/DQvpO0mdebzWI4VRSfrJWMyEMikxZPqCR8bFW4KZLK8Mb
VXAG6c75J/KuayQkjtDz/VETsgweyIG0tvzUNZlVS0NbrCd0DbS/+OCSVQY3b9KrfpqW5Ug4vQTI
uYmhvPEwVGW1We4JL44fH3eqF2m1yyMCS1t+6m8fadyl2z2mfvBiPvCnp0W6TjdsLNS3jLYeEJam
7oeF9Q+2zlFU5kfqRziPyQM5ObBdREzzZD7spF9lVlOmzCN1arubdynijjzfNDTXSrxlksTAAh5D
XuLE8bKEi1CBNFoi7qzGpLtoas5G9yd6v7EggbVEGhcTuN9zoJOdePviTZwR4JJegLJXh5tuFl6o
wWdSQ5TFcu01Q48fo5hmol+sCI9QsWi+wT3lLOokqkqLFGqf7y5IYJ8CAz9HspAZLIijzfKFgNQH
ZEewGGXGa1TqFXAppsJsFAg/jm5dynH6VQ3fcB2q8soLE8aa0QgBXh3lD/N+rgYB3MbCG6q/ynGF
PHignWeiQdAfyLH02i+hvyRPd/qV8dowMWvDpPrdfSHNDXTMZU+Kdn1DcSRiRi1E2upQe7rcEQ+X
rgMLATa0YkaUgZXz0tnuSEs9rWdaunpl0XZBcVVfqzRU1UjAa/y1FNMaFhLGh7oeJj6v8DT697li
NTMAMJPSmeiEkXhHVQ0w6cP2sTKPmTCThbYtz3Y7Fv4quN5M2jdEOGeflABtqJlsaH4BQ96oarwv
0iSDMgqmsIJdYWdYggz2520FVHpyM6qM4QNlCsTMh0bKJC9HEJ/bb9ZbFqiO2LOXO5RICvzLY1r3
f2GXveYuJMw8U6wwKzYjfENmPGB/Bvw00QY92tmow5nxD6My2xhy6AdhxP2PRMPOjvRePe8zDl3A
U7lolbWYkpJjyjkxvdk+kF8GcFh/Sei3/kM5wjcxwfV5g2cbMp/l0IMB3fKZSnO83JYbi/yjqE8M
PoBeqNioL5D+2BZexxy0fu1woonNC3REYsl07beOYPKLUiMxhQjd1pKmqcgrq5ZYX5M2MYvswoRi
qzut8M1SlsarsHvXoFE8FCZ95m+nlxmmn1zuov7eTiXtZUpho+AyUOncU9gz1Ph0BBMq5Yix4MqA
C1ryZRGRD4iSUrlYfIQi835J5SOkKDMWFTMnqKfHkrakkRQnzwn3O7lZiSdxVbMNfZwo0MGwKP/n
C9e25GRGnMxXYsqeqsPG7LbkVvF0M8Vua3i1hamt5zP4Wh17O+DyQaqLbnhB/4UIxc6j+yCTQCCI
Mbd98F9oy7tKw/U6ba5XH+OrUV0ZbI/GcVKqHPFgulXdt/tPA3+ySNJ79jhLehFs49BKkrAFu0jF
yOj6IiiQCr4ZaegfIU1sM9IZ+KyeU6kM/ea5zdPaANhio3O3zdxw6UkbslzMdxPHlDNb6tPISvna
jSSE/B6UHZ0MUl4oHdKO8XMURKBJqm4xyZEltM4ogC6rFPYjKK8HRErveJPD3MZoQVpbDhAG7VPj
nt3lmfODPbXvVwliDJyOEOGXLIeor24EB0WhzhUjj6QB5lUgKR35sPlmBwXtDYYzYub+qVxP4Tp+
XRh+eg7krTdFySPRpShN932pXDFbtm+nTnsxFemxMCXcUQEiV7dpxnuVmz5tCUIk/BLDYjNFUMOJ
d0f/GKnqgoA+9u962LH/JpAlhz11EynqS6mydu7XRcnJhp3Z4SARJRqsz+5pbT65p4GtXi8Kt9wd
Q8gUaR3QvxebFey6idFno75Ad9+q9whKzD2g5HTVhIge82oGHij4k7xkpHxIigxsdhhC6uhaBPK+
CabM01Nj+6alItdTdMZctrgEmPZkMFSDpuQCxaB2Xmsas7MXLYsbZWsuZTaowSUbnqQSWsQysRXD
+DHWTS5FTFBZ94mpVDhnik93uESr/5Gs6pkqc+zZpW18u0gJe8XdvoQ2Sgyd0UeihHWOmeQwqko/
MjfuSlmtkNuFXyUE5SrWQ8WYFwzSmBh00wH08OKfxCP2Mqjf0fk715nO+cHdaZapVj15dBg8NzZv
ivIAO/hQ29D8zPm0UPSgsObGoEoSYTG40vM6OAJvTzAHfdZZRbVpIBQCUbZ04fTEIcmfVcqG0XoH
YQsDWgNl4vBmMwkZSE6rZQn5eWKP7+4pvNHAYdSKg7rc/45hauofnX1qNyfvnsiZY2/6pbhgPxxu
+aHbQXwo4IfcTwA9n7L/Xzu8TWfLXXj/0pM0xvXElOEmYPZDA2wOYOeJ4fx8os7P5qIuHz/UdYoY
G9Hk39EpNt2Pbum6P/kqcKtYXgzKT6w85/jrecSM5gt47vx6Ii0H7Xr1o5rdWoHgxjPPZjNcraYk
6PsjyCe7K9Dz5Is7Y+O0CqZolD1huOsJtptyo+C1hbxvLucizvJxUhT0A2t1Cu1V7Ds55t0X+rns
1zXzuNF0sHxqqQ821dk6nxnyu4Dv6n5d7ya2gzP3sHxLCfCeQEAv6kektJ88ACxvro2WXtfxeyin
D8LnunGheQLxsoJUbxc3HsLahwfD4mdABbSALyAR10ynnxvYczjbrgLy138IHRwrkJJBvQEYkUT1
oG7AlVzPuYsipK6axQx5xwFX5Q3X4seEzzY9hO6sVXja+4+JLOaj0vryd+vZL+it9ndDTwZPCcV4
O5ODSOKM3pTBEtIv+QOKoWi+Ow9nGICZpBTjFJ+JZe3tQXr+Di6vFsbU2QrMblvAvZ95NCzL769I
mtejcTzOXr+1P09r5LQIhuq9L/dzoC3MI2Ob3Jh2hEMsmZv3EPm/BNA2kyrfs9rMUl2bSRy7pTt8
8KiH85nuVGxojr1RkC0TuMxA4ExCgTgO0OyBmicQ0Pe/VByretuf+ZENwsBvyg9ysuQQd6ZKBzQ4
FTjNPctxQPOUhlWrBx560kJPQRPLF3jBHFK6k9DbY9Bz5tawrxLXXrjduwwSNqQWDlsi+IXWmaQN
gYLmZ9y5kCtdkdgDBWGmW4eXJQk8Qwn7l5q/FsNdbFEziSWA7PddVLBXeTDqVOWWz4G42C9tJn8Y
/9+x80H9CiaVhOyyeGME1HTbEswUP2nRIy8lHA89/rvQbFlus3VHP4Vea2ldil7GCjMYppmsa1XN
VSq2BbRuJV5N5idtarJM57XIGnm4Iqq0zQq8V3gM2PQdI4fAxa8XhpXE+PHJ7LyUnLt5w+gZvQAQ
zlc6Kr204BgKs5lAzGPr4MWGtxiyu76+cXC2w4ZMaxgs8JTIFaQN6fuUHqkQKGYCbe2a6n4wfBZq
c5pYiExhuiP9UrmBiDx7+1hPI7pztR8AfHIJozpsDGoh9MWN5kho9vSZB58Cr+GNW/8EB893Mr6V
+MQFEDOsIFPkEKagm7rqWl3IVFfO/1WCe/yl4myKbSnOLf1dLg9QfjelujAAyTy6Rn9I0uG6/fP4
gtW/jRMyJoUA+9L9gpAK5i6BvdbTh7SA0rOc44XjBCjkOMJ1CmdOVRwtqoNS6OtP9WDTdL8cEX3i
oEh2W80UWviq9OQtZCwl20/W0ahGNlXs67fE/i9TrUevWUIGbYGEemG3edrO2SXZ2FV6PxRTFDOs
T/aZ3sttxz/6rEBOtwt7VEtLoeIKwC5M6udqoNSSEu557YCx3BpbPkuIvfUdKWQapDB0IJfeccu7
K1DgbQNqN7kgfZwiXqo6pmX9NyOCZD9mha8wSDb1OGx3OcDiQtU+ORzoZCE2OGOCpaq858zArU8B
2xozEz3aMcKerWG9sjHA12NbZ4os7au7bUHgVaHXtgw6NoV1JzTWkJgJ4bsdins+6f38cf1dScFw
bRaoH+wQpZOSKCzVixYBTCSwQh3nptjXl1F/hkWI/uPlIqPv6a4UjpuD4sINkJuBRWmeMrmfZbj9
lcgxBF5uS2xcKn5G+WXBI524dBGDzRtfQTQCRFKxMTIlZmWIvcFCtfwfVZihuxYzAsmsZWT6fDIp
6y23dkfjks/nUZJjxKlTye9c0x2WnxEiUVBt3iN1uEaJx4J5d7OWdW0jkapQuLOWeYwJIy4P5xOR
bt3GBxDzIJwKgXDR8tJ1CwHybssgBy7kXZz9cuLARWHQR/9/rnJE40Apta9NYXfXN30WCTl/82iu
EvkuP4FUMOn+ksoQTpcG7ROH0G8cF4OYOcg+oRpddh9oKoCOl5M8WTe8w0ZsJuKrCvniWGCrDSzb
vY3A6yxTtXnjnv3VlVP2/1CPWqPpQld54Ocmvx94lXMnQIAs9HoTkJh0QYbTHUhgvg1T/IXsYiip
xvawC7Lk3ISHOdeyeb+bsGPz2fgASUQD0cvV/oVOtRZZSuM1Ci+eSQyvwVU66fF7Hz2+wJH02RjC
xWfsyBytz4ZUSqnhbp0m/UilI8mSAbGj+Igh2T7YB7l/AceZjz05dsgsOgM+8sz/yxhgIFNgPYRa
A79UL19UjZn5/2irx3BZFbfz+zwdddJkkqDsRovUvHylu8lTAZCoIq0wItiYUDpAb/Ab4oUP0CLD
i7Vn8fDVwvYCoAKo9ecR3bFK9PA7UdDZ79nTFAJZkb237JoCzVaAHSOLSAcDo7sTCn8naXIEUIj0
ARDworuJ9ziAiarONCxI3q73/dRU1CARYznZZ2TTqhi+ylikOemDMjD63GQxJBqfZRzKcC4eMfMY
CTPejKOXqCKbElXq8cY/8JKg5I2csqDguZ3v4b3F6p6kqiTpklRgfJe5jBdkw89JjKjhfzuoBHxq
CTjUEMH1oVskfFy/84+xcHnlc8naKKX+iaMh2ZdpMMoO/BLdrnROJfioolk2hrKFurxvHcFxIYVn
6LHVUrYwIP3QzyQO/rTAAlNnXmLmJuGZWwG7v6a+xIxsO/xEfjEWC54gyxwL5oEEsDDtsEEHd+cI
CBdOHZHh9ZVWyXWXGdA3W/qEc+2tAYgFoZ9wrP1GnUBtehVA/o3UyZTUYpnR0YK1BbrHkWTZU1Lh
hd9mJuW9W3G7UicsQqzzBFOnunZ/PZviujPiSUg/pmDzS90tU2ICtUExVEmV8faupxgjS1AY5+k7
jG12irZIIMfNCR8t8g2qLYU2CUk5EMwdxZ0jD7v4pdCjZjPopasVment9BzuO3S9rlBElveeHaJS
lS17xWStPU1M5i9DgUjqH3KL7fmu+bccGYi7oadjXiUvnRqJ+lUSe3OqR6HtW4u8aTBCol1i5+dU
ne3ZxIIc6tcVwLk+OnfBl0HS+ua6s4/6ONkNC9apS3tp4P2tvIXMZDkgtsKWF4oHyX8u+JQMW4GG
P/xssmGk3BrI8eno4nbLZvHtEfQimq9OnQChCL4t0ZF0nWkC8uj7GZPoHmUJ1fgIuhLqdw04+GDg
7MoxT6VjdaBqwe7DgABO5tftiDmjRhD0SDQbQl+6tkH8IV9qXKypBxaCUqGyTP0cQR1VcerDsLNv
jce8ymXJ1t0zY8IeEGIzlzdBGi3AVSo7ezfSrUICpNydiSalZ/j7TZj5mkq0PH8Vcu00MCzKq4/n
UX6ilaWDTf8WMhQ5fdybl3jzdvq0Zv7eIVoCzPpzqTDIkR3qB3OU06cdIGIGAxbhZrsrvVF1jXvL
r0BkhwyJh8DS923pRt1UOQ1fT21swH2GmqSXJM33UqMmKVN950QAGdZCbUkZvg8hx4fHtbZ3CZsi
5YXR+M0rld0EaiR1x3/zJt6L5j5xfFNZvG2f0RyYPb7W/RJyoo7VyKZpQfpKLPado5ILbGQbz1/J
Cs8YSQNPdD2UfTkoTq6oyyzkmdeh5/rDREZhuYSrX79ss9+vRbQ94PHuy0h4apD6aFnRT1onrkSD
pJIjLnPLxbdFiPJeM8G34ywpk+bL5ZMs0+AYdiT7nxJoFVIAvmZ3byq5UYlt9x9uloMrMipeXmB9
zaEMHnTDDRsQi9fZ+1jgnDY0XFEHPCT6nCrDLlh3JELHDZ4mYaWFuTmzgxclgBzc+1FItMWkiIpd
Z5EWTjtKgCcjnt/qUZu4RLG6yjJGpiA3VUAvtp2NWk8HaYp7RnFPGiedqnhGMizDVhemrwd8pRXX
cGgD9a/Bo44rDyGU0nFpamS2k93pnEuj5tDhN9h9U8fYRrZF/xPHVRAd910oI2aOgsD7FXYVUpV1
yOAucCdTE1aJIAPPcf30QgdbYZMKxo3MewOghdyvjesaO8MNUqTOCBAqgtYvC3LsRg29PAn1Y48b
WXdvH2BZkU6Y3awJf4Pvs6I4uCnzdNxk6OaLZNP8oyaL5vg+o/p6eCYOqUsXfLtthzhohFHMLTSx
dD6kRQbNwF3tvvPeVeEAQ37USxufNztDgjvH0Fzl8LTb/tjZDTych0fmFzVeHJ9dKZVYwR8wEgMp
MJHsoirIOWDIBMo67qDnM/c+NBhiWN7wg7Gpr93o9WgJpGfQ45w6RmgqqyF0TQF8wuHFfVtoTrNU
dKq4cnwwcodY8Ya6e85HvA6yX46v5UoMQ0ILMX6udmpxhxeGdGIXrT6C/CPkun1fdl6tNzXk4KiG
yvfuKG2LZpkhDM0VIcSx1vXH7acSmCmZftuZlslYzWIcqepEF0fwgt2eV1IVD0CVObMVVyx3kXTl
Vx4ArZii831FwlFoIqbqmLOt4WUjoGGDTnDisz/TFxcoL2mrj3fE88hOXE4K0TaEOKaevkxAEVBk
l15sOZrB5OYSiHtOxcv3dfFNUP8DNEymxavfw4uDLLJBlnitNhJ8Rl0ig8J1JEh8tqXtGXhGh5Xy
pE5JX7bGtNPNEGLWBs5rhpE+bDA7UxoMQP98oLS3KTvHMPuVsM5eccA5uJ8H0z3Mim8ViH7pMO6P
jTCmPlqR2nSchB+7IAfhs8zAMtwxmu8F6fgtynLwjZI2cYp/kiQIzdlzz0qm9iCkZWz4LD2dnKzI
XfMhHwEjbADN/glI+nIBCGXGEByGS38Aem0MvHlf8rqhTzL13bOEY4rFbcyiEbbxR4hKGUblg9vW
ELtZZODA079kxO9otfSIMbTBi8gxrHxqASxZwHbQMcHDzh9+8y9yOuSEDn+b8kcCloQ2kNHz/3SX
rsO6r6OfLhiUoswdeQOZpDFLyFxvsjLwrNE9T1MNnCOxIffqjOooi2pSmom/1FLHUxpTEt/NvDbQ
yu84CIPXswIbnKwiArqs46e3bxekFIUUcOEaavdJ4cpcIakKjOenoR2ZIZvwUKAhRqSwLxTfgVRJ
a2dEB8dHD2yQwA5RwfQZ4trCKhmXZm16UEN4k+1WDUA4Sr0sy6qJ+wFyKwas4KqAoURXGYJpcZWv
SuxIjbq7ZNQoejkBBwilEJU4ZGJU6kQiIhWmFXOb/MsKgOczYn9C9xx+CBnWoSQQF8NIbLNVJ0IZ
okyHFrOgpBoCqISfbWqP/xC8C9ILX0UVWY3tO7L/gT8v4FQOw7sWwAUDLxipw6X7r8oYj60YPaia
onTkC21LSNHZ93VN9Nq0xFldGds6UwP/rSoCjGMVUcCHO/kef5PbOd9GLTepcpi68W8C174+94eV
6D7LjWJZX93bgbIEP29ey7MkGMbercn/Jlz8S4aDbfZvwogbEj3Mn94zr+Werzj6EeJ8yjD1ybEx
A4nUnZqlP1GN4WQ12/Mk3N6iHu4U54NrkmvX2oyvrgZHqJ09E85hhA7P1B4EJLDgS3Hz9DBZCvhP
ltokFyPUo4TY1P3ivc2s6J/ysjVcnn50it7+Lj7VoGdVJW0m4eWYjCwBWfc3SJSKWqU45GOymCGs
CxwbGWozQJNTn+ujHOV72HS8yHh8Ubz9kL3X4T7QU/OGxKHHCxUhvRZQLjve9/Q1K78ZCcMZ5x+D
eV7BUoiUqsBjqMZKUfdJCkOqDwyuqkfcyBwWTYtEGpcjm+b6s2N4vPPDGbfdWFhzSPNgIpJAC/33
oMsUkapySfDStG9WT5DB0PrgVyJYpL53ehcJBnHS5DQeeRUKOeF9OCjeDq+dudp8fSOVoX53Jk5a
EDOBAWHsYoOYQ7xDBrkZ6OWQYugl68y1mqTkxYTPkxuPxHedh+YZ5YJU5Bh+suV0ulfoHt2bwN1V
vI2DQ8DwRpx0IgfD1odNE16hi8ZwIEQWlvtRIVHiz6Vospu3Mx6dLaY2OqcztcdlNkQpDQTYW5se
S0Xek7FAhWqVWgxcx25EmJPX0Kxu+zJTeaCRWvpOjwCuQt4sjHgn6mT2G2xhPyyrD8C+ecQEUATO
/L170RIQDI8NQWnjdPIX0MWczLdt4oCb3lolgpepmjWUQB4VrN1dn+aTnQTN5I+aBfud5iAQ4Cms
LVxbvRebzkZIL2j+y27wMxb7/USBjSMXQVPAoTvJUCtslPC/BBUJJ17NO9BY8ZiFsSncic6XD8DD
rVJn/cESUbLwirtDOny4lfUXYdlHelYW4O/n/B8igXlQ+sU2DJLZTZeUpJNbNIxqv4E7GPpVGpWj
h9y+zE/qMK7BplHW0N6mlPrbJxHv61mrzW3k0XZdRWNFbMhO8c1OthG1RrVAng1eeYYkayoQMkJk
wmR2Rnrj4NExAUq+cb4VpeDJOkTs0j/KFv3nz9rncFk2erNEaB+ixo2UAuRY5ty2Q/m5F07FO1+R
ilRG/a0beHDU6WGrH1AY0wt9bmBagIvJ3m9+NHUru7XG35xT14OuIFUSCUaAB+5bD2UJUPdVAKst
QQ1Vg9sVnjrhM9kaf0yEoD9wG0e9nDFc8tQK4kAeUqNpKVYSNdaUSQ782eLRZ6G1u+MPrigjxoWY
DuXYNBN2x350LFApUSNiTrNc1YRyF9gJvhwltM8/QMoIOmLRR8EovVO6CuKbUT4whNHcP1sbs1eU
RVkimaRNFydQMY6RdMdFzXsex8Be+OQ5YSFNx8pTbYMoFwdnMbyLaD/e81XKc97Z2ZXSiI/zkf1O
OMbY/YJ4puY/jKDjX8XwwgRkSvdcl4Agl1UjCVk5ciYuD8R7DRB4zEwSytbthezBYCwe2dp9jDK/
Q92B8aI79gREcR8yKJ+02+Rt4YdEcvgne6mFqyBLUf8BHf2/7h10cmwVmxamt9of93pW1QOo8a7u
ESAGJP3RkG780iQssSes78+mIy0k+K2Sn7buNEjNhRG1gfIlpFPfbuRUlAIBt3MVRXfit4OtGeAq
NR6sxUCogDZWhp8Bqx/a+5MoD+aJBPycVljkOHCh6mNrKqVUBpYjAK0EpK19EPXTNX8G8uUhlzvn
yYbNfl1KFI7aWJ07iKyHXM0NfD12YIByiekE0RNhu86TJHSlkJxJVOwSCQMsIT74NDoj80+9h3yC
PE3FuT2YMHYzuQwnPUK9e/9vAx/pN/pHB9A7p/Ew7B9jcgQApfofrhoE8DdL+iDCn+9BJmDq6/vX
T/4zg62OfivpfkSoqXF5KPceEORkwK9kAiTho1Nem3dUt11Ebe03pU8j91yJd+U/YtA6Ek7pPmpb
lP0/eD87aGSdZ14j5gDSvhL7MuFCAB9ltywp1WcezYVOCEw+PmOnm8B60LseosxN4p/lKkbZHo3W
SHn5oMrcGtC31Bnz+GpOA60SvmN2LxnEhfpD7uKwj2RL2CcBwjlyX9x2TJmIKs7efiyyE0RUnEIZ
B6hIxZnvR9REC+CGecNNr7brLEwuWle4wA+G+RXHabetp8roaQiSY7rwnF8PEOxwnxFGKW5IPSHe
jOaFAr96eUwDd8QKy+/O4CbkKS71Dsdu95oNsPc9hIHSJuDxLHoXSVvk1BqZidP/WdgU16wskmfw
03kJ/fqcCQSQUcPr6bQdgnwpDVQIirgKR0dfvNldPdpkRLKKtJA91DymdND6zluTcsvcNBjA5yEm
Xq245yymh5YkpGTmNbc3QfUzVF4uKTTvoJeWiFvcw0wEYucFyVmdlCbjrnvAxMgakcy5Ze0hDRJC
r+kVATO7UA9Wdxvmx3YLqCGHlVfsMUv1eLCzpEzKAy3GwbrR58uQH/VRZjj2285JqrmzxvWJXWhQ
Fw/8MneBxEWYdyQLS+hBuDjFF3GAmMOFRFcHml1uFpR5KsWvpDT4qdEcvB9eoIIR2l/UhXJ4Qg+O
xPH7Zd3CXTlHVnCAbAHADXz+FyhwDqr1k5XeP5VxTHs80diL/kmZoQo8j4i/13kd8IWbwKctQ4di
7azJkCYpVORt5qWsf3jJ5/fD4GFZ+b+VRJHIO58tSnljrzVDnrhi2GrZGp8lSbiKsnQFYThARrU/
9WnA3Nw3iyQTcbKR/i9A1wbK2goKRg54Yf1n/YuNMnhF3NWzJeFNQ1wE0vZMaQb8l9XyhRqlj3zd
w68fPNZ3oNzEM7im4Ybz+XtsZdlfceKQcKt4xqd9yIiKB7Hm11vCsUmRusfi43XA8df8d65J0fNC
rGuM+7E/+khGI8hG5sh3d6VTw+BN5vn16yTYvDwUUcfSvZeV0WKkX+0y7K+1GQGOmMQlX2qOHS7T
6EsDw24DPFoM0CewwbMb/+2DEEw97a0HZ+pFauFs+XlniP883+n12bcvrbKT1OoUtT5HNo9XAdBX
8aKLsgfYfUTY2LJ1cUCwcXG7CLJrvgLrFkKiK99kQ6W3ikuzV2oFAammLLtO0I39oN61CTvGNE7A
qtzwP9p+v/OSDpgI2EviMGQloxCqb0xJ+XAxnVdm1TN/s6QcChKdwrs4KAEGCBCpgz4P7AKAZ00g
afB+bLd+zWnH7uEnq9FwssY6aE01TJRit130K2/sdo8zqu7LpsI9q1+p/3pFaXq+jKvjXMXplR9I
aPX1H5MHqJswRLGuAFtFpaFneTnwSjMS0xccgM7HLvDlV5uzMAep6RH0GxmFV9VAONAHYP6seD5V
cd3LP5RJJcx9qJ4CWtGM21ycsnz/nMdVuhK9yO2jQHSNZmfY2tMwc0NKiTLT/7oWzfnTtTaFmRxG
JqORQtWbOCTQbXp/JfOA/tiTs6GWC4SiY/hTzBZNKNr6syH7vhwRrbXAYKvXCxY9RwMk7/sTO6Vd
wsTHtkqymcrMOWxgJZdE+uXzHremsVpw4Le0WvZHlzfPe68cbx/AntU8QSf9Yp3Z0Uck0oWI7NmB
28ovzrrAGszRwy84kFXNks8KHiC3XX2+B6Oe/Cw/m+9bv7EhwNGm/bXjQNSyk2/WmCyI41QLw8au
Li01genbpmB0JUUpJqhHEGHLGtO0Dkh0EUv4UOiM8LmVPtHPT89hBzIkLptm841xv2V1FsisDJzx
tiZVc7dLvUmWkjnxlva3LxCs+RVVUcIo1y+qNRcHebGAy8ew9Gp7sBll8V/lj8jPxga1AAhoTM0y
XpdxxYhFXqy5tKBcBq2cRRgXL8/XoG/bokl6ONNWbkL6BfdlAQgq6VMWuHTNJXY+Zzdl6Xqbtygf
9bJUvf8kYUIJEzyeJD3KYTLiyK5EB63g3m+DCVU2D5VS1HNWyCft8qH7lPgKElZ+owc5CampG5/f
9tGR2//YwLL6BhSrqxkrU8q5PekHf0vPsxa1/7x9sdV0pbDtcdccvM7euWsLQQfbMt1/AzNOJo9B
JvUzFVIbc4H55hICoBjMLgqrtN2inFXY8EtHvhjAH0x00xVRnzvA46hamZM4I3A9a37yHuWl/+yB
rsQk/ueiObI8+0panGsG/4hpubFvCCCOp3ROa8KM/b3ecLM7wSTaYhzTHcnxM3PfzXfa968F44Tp
k4uHAFxy7C7j8cacY4yp36JuEKeWtEDU9/XHzQpdK8Tg8rJIC6ohtF0RNflYmjEdCToDzt7SA8yr
+SUkKXPZ6vItYQQg+QNXMcjpgZh0W5VYyh7467dotb8XDCNfuuk8XXLhLttlcO4JN6iue/I6KNcD
jk8rDKTpNtOQXXK1/LtGGRAGlTtpxcGnLq/pWtwB4eyU7KAy0gx6fzAK5PesgtQVfgJrvr/NGJd7
Ix5sgB2CM5UAhN8w6g21bHEpoWxVdfR1bBAKhf8KL9KL1Wz4eom2a82qOUR8rPpx1UwkAL3HIEoF
E5axCrkd99kJ1bnCt0KDCaPpBhRBSCi5itaIgNEFoBL7od3nFXsKsUaNBSTq9/MdJkcm/xcKSuPH
Rq1WQ6ZrET7HXPRHsSUMpL5joIchHuddd+MmL7+IOze165+BP6Wp48Tpg5nygtI9+Cv1FjIfCviA
HLSc76i1RgdbEexFIWaCamoT7Bh/uvvqlFapAYGPCKSoXz03QA86b4j+tqBmcWub7IMnLx8GCt6Y
oTlXI9b8Vj55zts0Zo1X+tEhWlcxQBnxTmfNFJ0SRjRNBsgoKyXdAdLH5fk5zf0lC5qfw0x2xidH
btwJUAyqD2V2uxqV/57x/sz+TFi4uPNAvfvZiQsWOZpthHFgq5q56iwRsLu+vDMdm17R96YlIqPO
zVVQXa4oD/tQWTCjhs/3/s2X0DV5ssQYCbgHC+qYEwf1NqCOXVe0KADQEwfLjx3mIsDQGfSoey4/
NC5R6NuvLGEmTdKjnajfl5pqq99TYwg4vJPe1S6WlHxss/1lz5MN4EVN8P3kwgQGkrgkiicqsov4
BfnwdSs+x/yjTa0jQWIgY1VJXCxAXdGxOkAm9BC1pIOq6EUxrSwQs/pBqV42QoCSr3zOTZVXG6t8
N1M8ofEJDXrNwPbPHfJ48xyqAiYYgNQoD3d7m4xyO1PKCiAx5VxRyr1Lf4bsEMdccUMyvy53SWsj
RFgSSdJJMKJolGwpeDv1akYsOcU/xC0SWYsfG3aV3iAVhuVtlyTSXA6kDPY+Cxz+EyNUUhxM7Mv0
t7ZNTlKh1SCTEzBl8PeTpXSxdOGiXgJRuAVvsCYDHfxVOXVfaUJVLVYGAO9RKTyOm0sXWJwKkHIF
CgDa1J2Grz6oMXL6GNN+gXZcbgRBMrxepYV+uaetuG8BXLmNGBbhuFy/8D/Yz6JYZSVct1jSWpTc
ioMZ1b2pG4U4jQjy1vOgMndts44wXBAhObdA5ZowzykJHmJn7hIbB6P9mBjAEs3gqK7PtY11TXk6
kWAINeyH4Uvb45Hx74BiCjYsqFzhphMmD2G/Gy0Fwjj98hI/FFeSwTvYa9Oxvr9Dd64ricp+4evT
43lbpTBUMjaaPz3g1aSAunHF5F4ixGghpN3RULApuzxh4R3FrPi0Hr1h4MMeREo2CRoeR1xrH4K6
zH9R/tMcdbseKB/UkvnU3bBLJ2+jAwU5myhtHLbZzrI/hpYDiolJWpq0J8SJWvO6aMTBFnpeYOtz
SA0YDtsPlH7GTyX4E2nLH/p8TeW6vPiab9OUAZF3U1MqyIsvy2br+40z3pibKC/mEVJDyPx8DlTN
DmqNhnUqnBhTqRahh2s2fkzSzaf5caz4WK3jGdXl+otc6y7HO/BuNMwi1NvQw9tNZ6ZlnYZVGyrQ
VAGpRpJVza6inkRt0z+1As5X1sN2AcwSHuTFFWarVkmlDLTQXFXkbLlMXtPRwQ1yoXPeATN3/pBZ
LexQ/OgxMBd+P1GpMS/BPueK2dHCO0uj/mwurjZXVfc4Re2b5PwznK128cFVFwmxiv6wwedKvpcP
OMNjnuvs4qsovS6msUr/Utgg+eWZSxGRT4vd/BmKf+FPDVeIX2zBJ6dVnE/SEt8aUB4DbSInsibP
tLOwRYDZWThJik+zor7k9e7e8aa+TX/jDmsbjNrOSADqRVyuOnqrjzstVlxMNl2fjZ7Cqbig7tQC
h2vfdFqHqZ9mUfER6eKuDCnnrvpaVVn6hw0lO776XjdPtgZjGdY6H4x1fCbAg/kk0LxdiskrVWar
M2Q5R0YZkZJWh5T2hbPL8rT5PfqRyiXBThPyb845t0hnzUGr8Oe+Zo1g6sbILazr5H60okSeBRcN
z7Tob+F/PQprHuS5V10HmjxypVGQcvBKV7lFmqtJ/N37JITJuA46/t3ApomynkOemCoQe7FhahN6
hY1I7J2Au8sGkQ9ykj+ynRLSt7GnIdbdihn4fCLF0edjEWuQvgFzYQAvm5+W2ZuogO+F1gLePZXz
t8V7eDhZd8/sAo9Ibbf3x6YMZuhlCrbgBGFl1tev3fTXzobCrhZGAORpBrbnowLZYgu6y/9bQaqG
1ODLzKwJyV27Y2/fE8WspMCogW+euVpb71G4FJnfwBfKnzAm5yub0HQUzMtyA17MuoYqG3XqbA2Z
C55AKv7JjtWLX3HElHskY8jPXg4Z/4EDpxGuSF9Sl2PPfdz869zvjztUFsdKffcl7upME2qoFs/p
0ZJVUFsm7l8bEHeRW2z4649RN7zIuo6zlI4oFnQiIE77bg2w4xdS4RPojsAcaTchlOB3KC+Zbv3c
Qds05fzXcDCJxYrIHzZS407BVoAO2cS3qqd7pS1bgkTxbJgiaaBTGhruE2WdBQsYGgDs7CWHhqiO
geXETkWuz8Fy+N9joQBPoY+pXWQWg77YvWre9pgLEjQYvfWR+TtF85scNoiTzRYupGGLlnaUgR5a
0CgWeKPbM8pKsmK8PhEEzOGiXaITTWotUVxjRyMNH+n54ewfW50rdcEvKylWfKBg8hpOU3jXMS66
HKuoXbIOxCVkDTZWnRHq+0I3BzgnCXOdXdybi09RBNAaAfnzJVfjlL8TJh4Y+XnaMkGTWvy8yMru
7gOyIJvn4p1u0WgM7SG8lmvF5l4h0EOXJhDUcdQowTrVj0zY73jxPdMJA/mbiNoKVXJDfuVCMzRe
4aEIVwGyoLXL/yh4FaG0I97KNrv/t5gy3Y0w51ymRTXshu3QEnE2L6bRImiu4+3QzxoXsxGYahaD
jR/XURpPa9xPRfBBNlpg0u3K3Kjv7/y7+51/iTA9dzFJudv9XYcYbTbY+AO8K/e3oWn0NrIyHDha
kI0s9l2M6DGPkSPhnsyzLP9iNiVn4nLIy1LJXJ+ux90xIuoUegdpcdGO0IdnPfJsszS1Uxaixl+3
Jpc0D+hu5ghhajfxP8JsMePHpiGjm2wfPXxNKofZ2kWLyGY7BNhSBtwL9GlHn8bQyxB9Ce6DIi4M
a7d1tcpxPA3D/GIF/g8eHcHkA9Q9KaCa9cO6J15BWao6uj7zqOG1wW4nf1ZFs79V3NOIenVtG+6A
ay3keROsTCU8eWftnoBYvp0NGFmNyrwIxJTNa0k679GL0xk8qY3lJg/PawXGNsM8R6CgUus9qciJ
/5YI/Wdl2U5KmIK7g9JrHiiSq7k1gohBPIGa2W0rcBGs07NS4DjUVFll6KPF2Hv88uL46lXOsb2N
BZCEIAeA7a/n5JDKoLDmQTjLHlsHxsewbn2guCYwIOMJwKH5DNp5XBAntkmZ0jjFKo3ssV0bkJC8
y5nKLOB320j04C8pHBCddoIfOGF1j5gSq+fwYbhgsTdvA3lj4ovGJ4/53j8mhe9yM/wG7faIJh5t
K8xPUELtT/5NMem+OL+d0qNJebdITbjFHWBthWEWp9c1UaMcM8aZFgkpVfrKFfsyZ6uO7ZV+arNo
e9E72Phy2O4uhkR2OekrRFaMV3vj+p95GSHJFj7g0O0uDjjZ5AmShbLPj60jRWSTaks8l7gHc9rR
l7GkVo74RLu/SqZNb/ubIoMLdZKTHHYNyTbVoSho9Gf0kjjwsBhP+7q0rLv86MPlYDiuChIJe7lr
cqVOWo2ZdO69T5PvgPQwdUYa8hscbzDm+D/WIbhMCRKrU13dZc5/JkNwCXmXveQws1b4NaZk+Hsy
7kHbBMNbjjvUyobwd/WjJuoOhjyeJ2k6b+wLOcqshBdFjc/J32vEKNgj8xsxw8QPRyNAgy+bl+qk
dql/6xG0dMe3mjdVswjrzDyNBI7em7EhLUj8K37eCJch7bArRLxv/GLJ65mWAygBPovRzpI8jD61
axHo+5nKtwFiCQSjKzR0TWw5Xb9OP2QdJHy5oOZ7oRtft9YPL2hVqZtWfdzBt3MN5WnpwYAmH2bx
oR5ZWkI6JbLRjOUnHj/VJ1L+85/owvK442O4Vtd3Si8YNbVA4hGn1JrGNCOMdu/dDiXy/iMaKamz
WBtsjRc29DBxsAX0/Zcwognn2R3nN0RcjmQ+HmmKtBK1X1G8xrmbNPxfUfNwQMitSun5xeS5AYvQ
wWnWKoEhNuCQk9DandEqiRT8x6psnQcsoLZN7tm00Smrc/hSvR6GbByBObi2OXHJkRccYcRiHA8w
0xQ35fSWl7u/w9mQVOeWbgqAXBBrDZZnf4n6Y1adFoCOtRVrv+a/Wv7oaaWkmjAUOicu9OdPY4JK
AK0y/SpBcMxQ/hAEZFrb/kj1qgS5hqQGduoSNFTGmUNyhkaoMBC3RDeCafGFb4Fj8Og2Po+bkjmQ
oNodVUQbaIf2tbELJfonrixc0tZueyOtQgv1M09/UKalkip8CzDXdGlMW7A/JtKclAaQ9DQy3zMV
N6FmZuyMDVp7agmXCQOpmhBgY7qypUGsHqqYcl3Lx4Ut+0sW0844rl5ZVudda1bYHqXI5sT5FiNw
nBL7SPHdXKqwy7qmddrc+TB75FxkqAgBC/xNBq61miMIy5uFPcfVP3S5tsIdFCqOQAzRG6n+P1+G
c+UZbV4kY+dpj3FbQmPO1JorOzc+lrG8e87nijV4HZX8OQp/pvRmLmwJ/6/vZYWe/7gc9l1+PXVA
hNcsutexYj3SlMjGp3YGYaYxzRKH/ff6rjVS2fWrkVjx4w6hch4HPYgwtLq1V+6Kz1+IS0RAWuIK
oF5bO/ec3y9BKKLnmdLkUN+wEde3Lq6ThXNbmpdL1xoCw2pLGgEmff50yuhF4IEwG9YzjH4xpYYS
kNgED+rt4vgjr7N5Skq9XWTECpRnTsVZY9FLlaRhQ1hIv23EsrhbHkBsv1eiDfnSocVIUXepv5+l
iel5+lPpoSu4qx+lskjocScU6kusOiQXBTsQI5LqOJp8vy+plSKuuxmutAKl0IXl8EgIebHZdCi4
nvY2QeW/UXVSNOqv4qlculhW2F1ADSZOl6qNzse5kibrIv3zt2YJ/0AdVYRR/dbz5+7Vy/I5K53x
wswZKDMgKa8RxkOWX55oymFy9WWxN0QqtgtGNcEKGR0IoKgKmuU7esrpK4sl2BzHZ1hLeJJJI7Bx
1wDm/9FrXPblpFiw3AnL2mYaS+RAteGgXdo8fjfCOen1Gsgk7PByq11C1MOnwGDHJbK0eLhuiQho
pVKqoEFLDZ/dkeWfEtD0Gs+D+wJpRRfngdRDoQRaoopfxdtJipjCOmW0ZDSBi4/7+UdVe20skXXR
qA5wQwbpKeYXGauTmJ4CsiwOjTwbwY8dbqBUd+8/ebdW7JkH/KkNvEpUc50rBqMhPLo+NDHinQGQ
vtTVW8AGgmoPypXyEAQ4rqyrUMOfV2TJ9/jtIby0855qG/1zk7nWauAwEtlDKsBXiN8r71oSvcIa
ruk8EZo4dYZGl+qQopPWPmLll4qUbIY4BoHt77h2uPfRv7YKc1ShLEPXX9ozvaRcyoldwkOLnxAN
6BFXuIG8U1svSaLqfeL0P9uREC33i69wH4SaE2N2xLnMtItbS48c+3zOFtq11nFxgVdJeHIVZKsc
kTm2CgnDF81yDRwfH150CMzube/u/W+Mk5oxe/LrZ4OPvhRoayVSb+eABsURROdV87vqZLBv0pm7
FaiOi9Dph5BDKgGdqgV+FkmLr7cBd2dFV+A6aYTGqVmzbH7WN2dtrf+6bGS5jAn7d/nenojtj5L8
n22jXQTZWy7ujAar4yP1mEUJcLM2zj8jqFZZI+OvJNBAqOQJk+eLrRiOmA7Xwn1Xc9fOkCF3v5tW
hADtDk4AAEkNgvWs3MCfEwoSqKW+rYPxHjJU/W4rqMOi4kZOBEZ32VdiytdVfl1DkKPdxZff+bR6
qKcKTjGqf6yQbSe6e9+6J5hg/R2xaZez0vZAGmeU3N1q/BARkn7TOlPtmq5zBikaYUfcsh/9RCuK
ASVlODVcnFOEhs/+6ljxsmQKoT428O1OuSKc5RBVkNU4+WEuFMxPFUmEcBMoQSVzVj1cLZF0XbP+
qpyHu/OQ/4SW8a1VZffOgVONMapIfThUCakFDYzkn6d6mcvdOiSGj+3bg1S/mPfM/8+VWnH9bGYk
To74wEygHvs9K4yo+x4DW3PL281QnbRyjrN5dC8zP8vyS8+xMrUU0ZuAPYfYt9seUhEy/aLTyus9
9CuvoEK/8w8SzFd1XU627FA4NNrbVaA1zA3/85ChSVfC9Dsk9nV757giV0QAWrGwyL//2fnFOHfu
yMpNEYOLi8eXPOp2jBkHYpqQnVoTosA/EE2nhOiMwFwM5dyGPFqgdufbfb3mMSTq9QF773hp8bjV
FYHiFdz5fOK6F1haKyrNJtmoJWdxpUebL+py/yjLexReDSeqBuAnGi5+mRLusThlx2C+wCmISHmU
1wNziJ1dWwcL4Zl+bNyMBFn8AlMLB0xhUDna/eXwiClDe67off+qCCIVpQCZH6FC5v0Zmr05zr3v
URDJlOCVLE6PP8mbT80Ypy0fayUBSG2c0HS2mkZQsXoUy8ScGlyifLQQNKp7KXWL7guaod7Z1j6p
EAkHOjnkcJRrSB6wKd0AIbiI+zVcCnE6nYuFQfJSYBl+X3BSMNYnBPZnbRfVT9aP6PZ+xsBe4/qW
2FZfBEL3S3CNnW/je2M5WOEWN15Jjhax7LITMnxUpis0EbwlesN3oXmxtqZ7gjlJ3fdrw52Bhxsf
lh3HQlQHUlCpAaPq+OElaFxbDycnsFFbR0n3u3otk47ge2Lp1mf68gIJa74e4fuwwaSMJzkBgL2x
fDA6W2AND7DBDHUkC5L2bXq8+37jLDlRY/PK0k4mSL28dRDtMSENZSuLadhbxUckl9ywFp6Y/Qzd
0K4dCTS+KUFCEBISY9SFP+64DYA+lLGF6dClki93EPmCuvpEgJIk9atAb5FdmxDKkWuZaIg+7XOu
VYDpglRLiBC8OuIhEjvq+f8WYT7RNZJrFcC2SIWnTPh/eMjdCbBKZaWyi/Spo7RXihCXQ8xJo3yp
dpAq4vUwsOGpOtTqE9SligGfVPHW76yVVOayLOjboJxNsefDUX2jhk8/1CxDiQsGNSFj5zFfIIlU
Q6wAUDT76v0Q23Ji4y4bFT4sJOAZ9nmaem+4hArQQ0fwy41He33FO8e2qjTar+802+mCxUA/faVa
aFHEg+hx1njaPEsBoSK4j9NcQxXZH8eQ/xDLce5dJawo/iv51REgug9QskKfiWXmnV4TF8g7J5aL
An4k5y/BZ3klGa0Lno/+rx9gGqjRTP646M+FpgbT4q0U4Bmnp2TQDmyQgxNe5ewJpll6ui1h/wQZ
Uu69zOXaKZQpbiL+t+VlJLpJ82pGmrSb7fa5V8jJ+IGjECYcXV9gq+B58Ag1Vc5UjW6jt8PN58tu
8qUu4PmWMaUVoK6id1GUwkQmkQl4SloQpljO4zMWCjFeKxKAgNf1X4qrAazP6IS3zcny3tABE6X7
8Ej77iP4AesY6OTIoD01MZK26enWl7znZqNQEb1UYfFpy4S73XTrA+xEpP6CMYJ+afbduqcabjRA
WTt+/hkQEq8UzK0J/oF0l1vhgqbybmVsYuq+P9tuAx8AeG1fMTdqW/o6grfPFbQ0qHl2+sbdx7/T
nl/iUQhkLBOrDpy/26OYxlynqQIhz3mThNpWr1vcWma4Ml8fvhCi/GZC63AQhhV2qgt0zcXEtKCp
jglw92vzL+NND2IS4fUVPzqm/9q/s60Xk1KJZZPls8yhGcPkA3H71x0e9084CtaovmYKDMSdp/jc
IMA8QjNiyz3IbxtRqs7QUT2MCox9v2CCAUmQB98R7IKpVnYkDGWpaucRSYpzKsc7WwOm6JwT0E2X
g1Fm0U4BbiOjrKASkgkelDBedFc6nw9PFl14eX0gbWp3V66E6mHeXavPD/Szphb2nZeXfU7nHZXq
zN2NrRUZD96Au9X2y8MNu0MoY7FJTfFVBam494k1GVU5uQTfX8msoQgxmfFOLSiUoBCO4HHzILrm
ivAr18Mcmx7wC+uZmb9FOP6/Ox8SuZ3BKXT8aGur0QhCBXdlI/zjLmorHJURJsdPNVjRN1/gsXwU
nVS9ZH4txsI3FKAfpozHL7rzsuLxXwGkaeUJiMfB4mxi5J781GEUpqlUYNwAfAPke4EK5ShEoGsS
y5YMtW2A0p9swHKUFaZbe4bdJ/RzDDglyixzWijegX0nimPMVTCxJtJEsTMZckO8hLNsTQ/Hpsjo
4KtyfCWIb2Db15VKFlHXiSx4vzLO5Zb0zMjcHl1iV05VVs8v7gx/+7gsl0Jz+KGy6kztKfGxRciC
sUqQK/Q8SseSmN7tXn3RG1f7rYP8dHt1bBkTv8mZ7RznyhrxH7lJv8WLHwAuX+WuCgJpk7l+25gI
mk2iesRxfOgxJStK8yc/et7S/DdCW+6xGTcMIfXo5NtZq5+zfLIzzbNATbjg78zJiiYSOrix5HM3
KJvWmKB/aqXTACSiwo0eREfu48ayI2F7EKnD+rqWoex7gWhvZnel5jC5vlqYIGdePMpvIvZSAaps
bqJTv5tNA4pKDPUn22EmgrqU+ZufCkZCPIUlI/O+t5vOtkneWkvq2Naq2sKjXQY/Poz/BJ7hf03L
cjcuNDS+qyrypOqDt6vDIMNk3630eRunwxMnwroL8s+g5OkNK9IXeDGQpHIiJDNhH8yHhpHPKyiK
e60Au6mleYJLSxNgAED1E4qOYPouh+ir9yYFsVF3x+GRmxTY2eRFLPd9XfFx45+8hN6G+iW61ArL
zB1a1+Q6lmKHKHzZ+XVUeG86ZJG37FPT3rLZELGGWGsCr5zXQZPVcAYGUssh4s8rBqoUIbOUIh/O
D9kQ8gjcMPvJblFlpoA8NYzwJRP3mt+r8y09zvbrlsQjev0H2e7rP2dM//yd6s8aSfwiqafK/LZJ
RyD1y1kwH1Sxr3Zd0mP21fDVCFMb8BDyQIKbdKb6HTdl2KTmPg2l4yBSidJcvnGaHP3K7bcdPG8m
GmA86EtSEUPoh5bX10hr9tKbn7IahbHK5UvVePK2gzvDtA6PJq4lRiQl82LR6UsfvVNMoGQz197U
qYbhkHj27Pe3TogY5d/0LngPe+M5Q8DiPWbWduiyOeUtLUrX7VYuy3WwSRW/vPL2ZSWXBxXtnAbN
jy81lx3lcq6kmvdXv0zR9D1tQSnPhlnD35RcrYuwQ9qCsKyPAGEAi2J+o+1PjQvJeuGQTYUT26It
JgzEn5K2oQhOdUaqIU0QbdHgitPR4wJfW/H8bYPHY8WGo6g72V32qHq96VZsTE/arMj7lu31y8hi
jIVdBvEzTF0jhOWlhydoXc5FRZaaPC9qmxMzJBhesUrKMZXtwuM/rSe5C2k1DAq7Tgd2/5O0lm9n
gRIZmXLx/46lbddFBesAwmVExn2p8WfKFwfFb2PJ7LHHq+lC+CpYfiyFm2wp6yFEH/4T3APQV645
xDRMv+ReQQKCG9dXstxKMsrTaDSuVG0iU0xV5vkNuRFmNQSAcMpS1NcOxs5y5a032M+tSoqAYdCS
4eoF3y6H6Dg7R1zWX77y/qVsEvh8pIYAO3+RQjflSUbUHE725f4CPrQZLb7MQEOHyIVfWEEoB7gf
Jcznot6bTbsPgY7WUuv8sdqIQjHcL92NsW0IqqzgImealorujE/qZSvqwUWp8t5tN7ri361QgXql
IuQ2dQxLB+tlt1Sb6/XbnyA3RoHfKMliDlqo4JEVMQ8aPf/SYQRSaI4P/B9d/jGDqtxsOImPOFyz
dqtKGfOJP6Vvo3JgDOwZme/UlI6H01cny6i4qrHxaSeppMxtlM1SQDGcIY35/68oNKxwEpvL39vq
umVus4YtZkbhRdUxisSObtsOtWdY+xw5IRmS6kkycSKkXOAL6+5s2hEQgPGmcCx8DDf7DEoiWnhg
hV6gZ1WA9cWdEKSSaW8DKY1sVBbfkCdxrp3Wqaj6G9MdJdFIuRMAtXsXJE9RR49F3+oy88cvJ5J2
Deu1oHWcH3Eb3F3OS4Tmajwz1Vr8lIYPgC0r4B19Gs7J8wCaYRYPAbSMKYIjrwh8tM6IW43CTZVJ
Rjwrr/gj3xE8qAyn2NL7zFwx3TE0Ws8/K5wYUvAhtGtC5DVu1hC6EImMPnEYUKoIT30T5gCnaV3p
ovNsknjweudTFBGW92KzTiq10N25VXcv8xW3sxjSOqpl72iroG6lIg0IbIf4axilB9jZYoeF23r6
7+8kNxvBuFVy0a53xeBRydjRHO19WamH2bCN9E5UuaKAjsZJabSZ2jwq7BFvnNIty9tBDs+aAlRS
D/1Yf3KpqLBcH1Gc9uk9hJqJA2lRFU5YeRE20x7mrS6DRaFEB3Wliaed7TPjlimTV2eVLv5mHqLz
Gz7j7D0jBLHTG/2yQQmE6jSVO+HORtx93xZSIQgvN+ylIaN6b2PcpmWEgy3H6szUdrKzzfqiGeb7
p1S7ClkoMrwD3ZM8f0OCuvO1EgraB4d+SaN9nkW/uD/a01K0GoutiYTvBKB0B/dvrpRWOLIZ81ao
hj0D7nOFYBOBwa5kFG9oEyyliIJ1IGfZl25aQhLpe/IZOlnCzeTmB1BQta8YOU8lGS2lLDDrt1UG
nj7kbn6lu7WfHuz44L48ZqHGVI93iVDBMtgjcfgbREKBN5RmtTRtYZMlSKm91A3eW+Dk8ar8wIEq
ovqcl1UBfWpvzf3E06U+tDckMfOk5hz5kP3wwHnEZnzvk/Yw5G1pjknzGGYpI71JeT2jfOpU+CiQ
egZsCHSJec/tpbDjmMi3WGfxV62mXjtsDuDtxKrZABY1vbkeyOpLxtFGeJ4Jhv52lnyXuVTnKgZ5
TPf15P/QXZkAG2oisN096T1jZzNq9aAbqA8OmoZq1n1Wul6XCj4UeQUt1sFktI+kgf9fbWoM3ejP
NY39XSaQv/qcdmghbjNCfX7cF6qPvjnvqKkCV6DoaFsu2gXWu8fX/V4nC0waj8ZrEw7sUir0ynMD
afmBJc/0V01BB6o8Ym7jBVLB8eiQw4g54CSRUgxKn0YYFzkF5VsYdZQphAtllG2FZPebHcx7FWv1
rk3FoouLW3GJm66txcongNYaZMo+f95DiCSxV5gxdOFQ2GNizqL80pS3zchm+ZmRMrm7vjcm8CX2
m4NX5IeGldjM/8dAsNMOpDvh1AlMMDXda8/t7SQBtmOoZlDV1g59ObPluHAzthKOdpAGDYRij60q
0vh/exGhmSO9chPrdIZewplb49M4rbhFrt9oVDztSogfBqCwvrL8AcYVxp79WzKmFzPtjvNvM8RA
SuPLeqNB5MgZA8ft1uXaqj9bVTi6VBID0tavs/H9pDU4ctrdiJqY8YPo8LcbBH0nqqhEvT4JMaM4
ghQbnv2Boo1QjG6Yn2Ev2uL34Q21jqdCLvZPAgDx56pxps0auC5Zne8EphXtsAvMuMLnGXTT5OuW
smwQ1skxAcTP7y441EgtYA13jBfNACx5QhbrhUuxj6os5KolQqIi5Hm7/J8oOi7zTRAzuNDmpwF3
Y2/HBwvy+kkpUTMUBEj5oqA8cl2ze/YLFZw76rXRN04END1FDZAnFIC5ndBTFQpSZSNzGwkLgoZ0
m9+YTUqzkFB31rF/WoWnECtLJNzhYJaXfmtPy3HWgAo5yyuJYsy/fgQVG9r1Mpp7Rq1mhl+Ht/ud
Lc166C+ueNXjXitFp7GMgTDQCDQEhMNIrWor5HMiWyW5x7LY40CAUhNpDcjDtJRkVwkTTQ7obVQx
siZwKxwN9X/c6OzmfHv9u8pEl+tKT6x+7k7oo73zT5jNCjln7P3a/RvZHSFPGBM6rqo341OQRl7M
AXFcIxb/jbu4vCqubP6ztbbJBqqHER5TTEv+6htQBvMswmB810kdseJl74RMYZ+Sw+/3owEO7D0/
E4gM7ikgJuVjel8tLc6NeI1G9ksm67x+38AF3pXmXHO3R7/4UPk7mQkQoFsjJb+CJVMDiNtab4Zz
W/U81pQwcTLB1tql3AZNXgi88NgQaceCeLLEx+weBzvBFPHPdnd+CXkC4yIlfmJTFuFJ7mpGsU/e
Tds4j4R7CYH0aeOfGgHf6j9iHO5018TDONZB+kuyE1p7fP/k+WbiSo6SNf4E8E4BY61yWHA7sQR1
7CvKbLVmt6d8cM5vBNUn15UjCjHaNjEpNBsfQoNsc9yasBrvF8mY41y4mF3XYCEBJuIkGufAjGqe
LoMJYTD4LOMjEMS/3eD3fathx8BZ2wqcWHKgaLcge4QGPVCGFb34/15rrSGQ8rNIsoFBW+Qejcld
CGCFJ7aTm9Yw2csr12VFJ754iZpcUAM/EyFirb/ThbQDmdN+SKA2spJfpTTgiLpsw2Kv6P1ez8gl
9mxDSlHgo3YZD1BqEDW1gko1cAdH2MW4N94OwLNmHjxtNnrcdyhB+B/Fpjh6zWE7dNOvF5j4Ccw9
pPssOVabrAcSfNmxx6ppQMnyikWP45LEw5BNHQv5qqci++Ka/hFsYNlv70ZcSkJXiYRiNqnE6ca7
ndhtJX3M9vELs7Udy3pnPQUKWvhmzxAFxFqSHSUYvxxoanCPdyRc9BgZ95vr0ALlRUmh2hZbgGTC
w/NSBLX3Qi+gdDhZ8lfxIUr68GjYldS2j1MNbepdTrrE+MBRNA3Jc9VCGMqYJFLI6hPCUGEvi69V
CIzIBvQs3VOFKJMj5RQqEbuPVX7+cm6IMsdE9Xqbbh5jFTMGgV1+Qb/e+nLIYXP0MQvIOrusXS++
qgy89l9Vh2+sfxsK7galWm2X3tX/+f7SuLPVGr7vYWB9on02aQlXI1Fc1GwnIEfe8HAG9oGs0Ulv
ksIhp2oAnOyOLL46QYBUHSrn4twW9MlMGUzzDvb/Bu2tSLZaZR8zF3SM0KQW7hH35eHawsZdStAI
iOe+oGRtj/RVltHlLB5jugUoayFes2QFJYxjZTydSmc4vmo5ai1fcqzv6HWetIhZDymWe0XNCNqd
/QNc5x6aJeq0xbRIDUX6qjuQji1DTHjnsCfAGXG2EDuJ1czMhXVsppZ0+Axa4B7Iq36xvvcXTIqf
GSWc6QRitcqEt+Er/D2pE5sztcEXo+Xnn2Zm5+cNdWLza9k6seFgsfUziSfSVnNSsnt+5ZSUlSQG
khCP+1Rlz/y+fTajdJxY3bYHKrPFtp4JQEmsCCUf2fcUJnEf3nt8ULECeEcqgkkkncWvNy2mncvn
EAv09NiFrlR3eoEp9dpGf4VJvbgF3LN276OxvZ+NhAjvj5aL6F8fMWCZSNacUv+9ZAaS5uTQS97/
z74JV4xLjRIQRVWLlGpu0+NUGGFrxqNS3qnB5a0VhOhweQ055CRVa4IWBqUvqAPd173Mw6Eamamg
MMJewm+re/ppZBR+A6fSHT32jTjk8ZFaISNKDz+W3hsQBonNAKKwduDoOVcNETIhA73HT2gNytQX
8sGSdsEylhM2YuOu/odJf1tFYfqFnmTqYr9+8zUHOSbibFijHTB1omkbFSIrSHaSdsxW1YJItMd5
ypAl7MhrryKWzLplcrP+T71Hn5EGa6Dyl6iA8kxsD/jaCbbs3x0e3O9RdhN4J3++DrcUyRcBNDCt
Bqwg+XgqwEDf2bU+nLJLT1EUFDwPtE1ZKMnG5YcQflRuEGtz6o72Y/Efr+aXP7WkWDU0DOjmPIuX
NDr2gCl8LfPT3i3ohrQ8Xs7GfT0ELli9IcoR4S008DuAYhMH8i3EXL83pe8hMkYOvh6uPOAUVV9Z
lQGTc6wTJqygEatT4HEeSHO21aZaETjIoMQL81H3QM+FTOMQJMrDYlZNJBOXCd5cS9t/yIs4mLnj
K/US/y3GOVrfnY5EYnxjqqQfCOu8u5MXSHJh0IBiFN2Nj8MVDYqRjiD/LYvkYz3yvm2IiiKxMEd5
VG8ln3vP1F28tfpX4bMvK1T+RkYJHq3meIQmNLbOhckT4cvqbbJbIC92D7Jn7uOWGsRveLgRgEKc
tLxzWSdtuAuLIAQDBDPy/hEqhNzxU0YO40We5y3El2dgrjGlgtLmFAus6VlkbMdt0zGQbNUw/bs2
HnDkc40xJAG7yS+51tMfHicyH2w13QQwUiQ7KmexW5JNYfakLjtThiGSIwv009fzvTBvKaSwSQBg
EHnnncK9Id6fgsSnkV5nMTWerG9CQEtWo8oBYcE/GcNxnpYLZ46q9Kf1LtLskTUgg9f968DAyQds
qsEj6p23J+TMC/WhYRY3HBaCSoVtG7qHuR4F27N/JVIExBRhrQAbgKsr1wAcm0hbvqfjl5r4cmny
auNsABs+/oyuy1HktIjjGUC4W7norZxZZJZRvkBhv6BWqTYNs7T1yhHbN85NWIe2o2IIAOR1X02j
QbuzRiCmhGYsXxutewPf+PNMYkc+hckqO/91Qd9Yk4fGxCZfSvU0jQHaNtjAe1BYwcizHlY6UvHe
0X3aFTrqglyQkaIVArmkmJOWD5Ucq1imWSWQbOmEgllSlEMGr5YAGGJOuv9C6fQ3uRKpT4mhJFX/
qrnGBWBFY8yH4AxgJa+pkz6aodTWaOGFj+Y1emUSgXHgERm3vAtQnaaOYcQx4+PTz4UmEgJ363NK
WoQ3tmb8kVyGg20n+TaAOZqa8jwIf9EK0ZpeYhZ9LZ0WAi3CF3t5G3ZHNw5xjoNIJf0aA8kgmTCB
F5zPU6lNvVIomjIsJ6mczby/uG+XvhClqx8LqMe8HvlnrZttnOyDyLwdyCad1YCT4uuN6BBM55U7
VNLgWuSgxjrMFUizLYPAi1wuANfcLwcy9aNji1N7B70QVtI2Jg6jbUpq4lfP4/Ct82C13yvbayxI
wNizk4M2fah8NJTj2n/qoI7yeaLEaylBYtOVkp5ZzjLaCxo/BD6elsRaOyfkR+yUMM7YXO3+5dvE
zcgVoG8SvFOvEw2LYHf6E6sZHDzmIA8r6l8r42lwjVqGYKU71A+y6ORDGZ2PGnGlFBm/a7RuKKbk
kihBZfhxssZZ6MyVlUm9Rdg9Ukj4Sgkd+gPW8U+rqmOYth/tvgVKT5B9C+Co4aaf5LxZi7HCPswN
OUX9HcWJ2wDYuKGOlhQaf1yAcKdWxVHL27qAAd3MoRg/R2LKItDVMpEpo/ewh8MX/LoQMN0CPdTm
p4Tx/WvLQj2kF2gTWqAG3ermAfODc9s4Hxecvkfccqnc7RhKiLFyAVUcIZuNegRcGe4sAjtZ9NDe
rG3BpVTYTk5niPS7vRwKC+1i1ZFdRi9xR5jOfoVo/lrEYp2gGYkR+4pIGHp3fDlmM/NT6942N0fe
mrM/NKAmZkwH+RY9m2nyve4nzCpysOcTGKvVNfzjc/DhXZHs/oRW3taSaAgnPfYGImyJerfFHeO6
pdSklkEoHYo+DzBxTpG7lNfRS8e1gS9ntuL1e01A7YKxajKS/9i2oeeMepVd7xhe6g4HZ/T1bY7+
UptH/rfS3GIgLuM3pC7sms1I2Z8kcJs8giC9ZIVC23+mUNM8MstVCz6hr8FRGrqHvi2N5AJ9Lg7H
WpTqku7ULhpEForols+hDwb52+hOw3/v5q5K96Yhkdv0Domj6Mc3eBwm+qqP6qljEXowAOVI6v7B
mwt0mZkWKuXPGiINLI/WEa44M2ob3V3IT3gITxmpYCSjW0kUbmlANStHqGd0I48H0mvyj05wWrNE
YD979R1RY23dSR7E2tcvIdxsLKnbAYG8iopyrFOK2Ok7+XyneFy/oCGtXckL3KmGIUmmEt5vIbYd
RGDRY/EAybAZ9m7Lj1JSpyGigTfCVIwuA/0yNDb2W/qWwwAjrRbb31JbPJC0n55SYbQbWYBX3PvL
7W2t4e5QN7oc7C9HX8yBWx40sls+dwO5TQbEELMcBiqWXL6lj0ls6N51uDtD/9O4bU/8shiItm+r
e/S3iG5apl2guv+5094nUQFxkQGk/hvN4giGUaOjtXJSJJwjDvrOuV2gjjYJDcfWbpXItsap9MwX
RF203NUlEVKWzW0uDlU/9vyvrhah/8Hh9HAnWZOCeEnzHuI23TIln0C5MVrcsJmQ98nWj72pgGWK
zoOrE9itdaRFKpXcm3VPwrhgVJ/vGShE1CHgHVp458XsIRp8lRJ8yl6ZbMniJk0aUrD+ATA0I38v
amiwDYQRYIdV5QvwhUI2uG/px+lVA+Ha0V2ezi30PGgS+m6tfzZBcrh6ccM0YOrm0/0T8l7UzRiR
hGbYyi5bHXU8/4kFGlGeDIRU0fsEUX9CLx72yzg8Ziq2M7u5x6xbvLBWg99FRXm6AhGF2oJxfz/V
MEYxe6QPmipA0/s/6QZfDdHD8kdr67uah7kwQOPv3NkgmfbMbt4raBz5wre4dQZSyZr4eh6Ui0Mi
ojyeEkxZYbosx30RAX+RgU20SaPVewKr42R/wQiMToGHwKmMw3qiad7Evsqs5BWbjGubdVu6shch
5Y7uyKcQfDNPW10FbhoAsbYNmQ6zdH8EMNgY5X8tnngh06zJj7/O+Kg+iLQPAuPQIat7KB+Gkqvf
88SnKtAGZw8WFjK+LgjtuhI5PDOQvYAcHt2PtjZm0/mf+CPbhlIdHWyi0NvqIrKi7bzajYT0Gi6P
pB+wuQaNAHrrPKoC/ytGI0C0o1hnlss9KQRTJ0IgoDXtQ3eUZFHBQHGgwBsPLOMgRde8SifsnVzx
gnklG5C1/0xdtzCUFRlTKqOFBo4tZ9VDJJq+01FViF0A3w0EEhhAqDMVKYxEamFoWOGCSH5QusOt
onSpx5p8PX+MJVTNXTr28DOX9MfK7fJ34jZzOqxEZrkoUKCCLZMn104QwxqDjAVhJolNfazDp4Ce
hPhplaj6pyNhaO8YfTWpbR73iTv5ZTSDTJEYWwFzUIdZ1BWB374t7l2LfMCmF4hoNwTdFMQnqoSp
QKdXEHl7nJzSJc9vy5mx/vW/bhsmOjmOD8NONHG3Q4H2TwDBffMiy2S38lcrEf3wD6bvFoV/EDDI
lYxFEc7Mej9wkgvUpuwKXQz+zFhz+chExnGORWrkIocJeE9L0ebc1h6jBDkWfceCAyk0TScICLip
5SIwsgTD1Z12nehhhSToHyPJKqhcU3A14zK0tbRG9tP/EfeDGQmhVcdhGBhZHzdxS9ccJzmC7/9d
0GPIg5YpkeewOqUYoUqpovd8MWw1QV5cpFsptm2eShDPPqF3m2zlIfHXDYPzTbg8UupHqbIEDXKo
GpqdSPg+PUzwOSObsdkRWP583O/OpKqYnxgwzRcwWIIN78PUFMNDRe2sA0Yo8kqoFilginn9vBZu
eWPEsDV0gWGh94QO3FdBBHpN3QO7fs9BAT0Yq8ftS/J0vT797SYL2s5pl8rKAh1cpnK0mC9jtFwl
3AJUfTX/buVAt1101sMqHZAhL4L3H4cq9m0uyuRo+UPrVQaGcl81+SwZUEhyJhHj0cGxoum3Sku9
MWQgTxnq0FJ6aH98hx8wNOdURULJqJXc+koXGeK2ek5OKT1DsJ1G6zt4jhHETfCJojtzwAfiAiRY
VwBetHS47tRSIMvt39nHEod4aum3fHbHWQoaorgwQDToCkceS47Lfht2NECEAQYWPGKbdI6pCDkM
Le2b2Csl5Reqa10a8pX8Vwf37S7URLMlVIzTgw5BFoBk0AOn0q8vidMHDMtnLIVzPlnI2yx/vsGL
Qzqj6THCZpUXeiHWRAlbDc39us72JnW6409RlDFAYhYKqIdC9L2gYeutT2q4u6J+mM2bfoJ4nomC
lVUh3UZBjVncQeXLog5tg7HODb+ll6uRi6HBJkku4zx4oyhLkkAIqosWjuKX7//zyrAREhTS4c2O
jrx2nIpc/cBywyRfY3gmaWGhe9+one4N2BGDRRjvib+NtKnSsOaG+xD2MV1uRKULZSHrZzhVFLPA
XC1dXgOzy8jxB1hhcUq7z35ld5AJB7b0NuUDHdRs0YndB9VOiDCYfvFLEbgewsL/aJM7aIpuodNS
ShCGxqOluHbzs7uln3uYiUV3mFkzoCc/Z13CA3we6r04UW7bTDPDQ4OtMC192syHP1oo/va13hf6
ngdBcnolVbXj+hnXUyrV8xBxIRtK8BSwCt49Dk2uwecyhh8DRquhSNLbiI+Z7oHoW628+j/SJF14
RWMyM0Nvfv/yvqI6CkwPa5ohPUU3/7UCdqMlVVqo7w3i5pWxpW0telylVAoTECTlJL+XR0WW2cYK
hnHV7og+FqvW+tUNUhzkqF/HVxURbAYsKLNQ8x+3umsd0cS0us8PazUluJ+ELhL0ITU6aBRKA7RK
deNnj2cd0X5XyACBSRJZYgNsLfS9Go5DY4ykje75CD0ZddoqC+vvOgTf4RLPYh2lWV/pZBJlP2c/
+i8pzlC9VnRBR5KERdsnV7+R8llKV91j6F1+9Sd50fFiTfb/unQCcPr9W+9rgaQUWKWj39qI5QdE
XXT5CW4OgUEPqMMcoo6t3rLMfk4CMM4ZaXiE0dMITslae5d83Fo4T+RbJkLK4nHccb+Iwu6USftx
Tv/6ABYgpyTwWZ0Lrzb2Vrdgay5GgWyx0KOkMYs3JBcPvqbfQJ4C9YEM4K7JMn2pgru8EiN8HSkU
peCWmTrWRp69sWI8qQutyLP9Bbtf4lFnWfc8e+q1Wx6d2WJaVvs0K9Gne8Wa9RiX48Zj6J41qvRl
VzaBrgkgckfSDFUAU+dCDASzg3uyMejNLXIrT981pTAvAaYaHLwsYCYg9nllyO8CVwNYQxxH4ehG
hkwBbfcFIL8jJmsOK6itXVtcCaJIKsoowffJvCw6Q0tuclV7drsp826Ph5QLsBZuxQpNCPsc2pFw
ngHXxEWFsh457mJ2I5IV6Y6Cf5Xk5nWMHkcGN0f+98eFsQLDjjyGofF0RENIR+LYgzrjxVNxh32v
fFiY40fmk9D6+9mHmjy4SyQtbc1Hw4AkimEheX+T/JaXZnjL/fHZ35NUq/RUKcTZ1x1oedoAinx+
T79ABYDYLTw/moetpYp7bJefSgXr/VR7pphJyvucHjR4G/kqyHN42PaEtFgsuZZvNaHfTE7hkiKA
1rv2PjMutTCMdMg8O1n/B/3MvKPxplGrtZb6c8q/6GB0Egb0pjrzgNloM/qyf4NjxBuZYI5wWGN9
Pqb/25NQNQ39qczJQBQ/Jeg4DoIwSFiXYN3+fNBjWywWprmUGOkP8CNa4l298DmMGKl6JOX5HQ/S
gxnNW52+U6GWGiNJvcTmbf7WaTKyMqmca3zRrEGiv90VaUyXAduHs1L7RMONh5vWiIlOXv0l2ldX
MifP910JkpM87KZocNUeHPiiJ+t59WnKWSDi0kG3wHmhltU8USF1BkEZNFiygZTYJyDqLF5czsKB
JAxpUmIIHo6Bfr4C3gQ4gP6WHZFf20sfNkABfeOt+iq8tJ1sz/xfGZ0HrLCxDKBBc/cVHXYPhDag
0WLUHEjs89WCwIUihPlZ8r3SygC7T33AB5+t81m0zOU9gOx/6uo2kCiyR8X5r5uklmE4ycalBRNA
tetU/rxr+BnKidL6/vqUnh9Q4aabs8ifJMq78Zzj3uzyQfThcz+RJ21hstetsq+vyhjhb4VY43nD
JL6lQMJvNHyoTIZt5HKu5kuf3T7EY0KKhD5F1XrKrS1eilKY7LN4zdSYFN86OfaHxneMPqT8KMVa
C1j85g0JH0Pgfm+pHVCW1OEicVGNLIpGAffT9dtnbGUaNKjwBMWvgZQFOkCLzDy7VRg0HCIolfFl
Bbg8MaHT1Gcs7lkLw+qbyGZBuWBOpAa4YqeXIZBIAIsLKPuj539Rjhut2hi+I4fpyor5ykf+ChsN
NvHo5zKffzkNQsROM0H98/yauwkFCOU1lZwzQofLFQH4orWK6jdCY9QplBNmHJ+5s83JR6/iXGjS
N2/d3FhHK0ZUtJDM2ltojiQ1d8Dzw6IC+jBncKDfhwAnyaDVOvUB6d51ctGdDUyR02C7qU3GR9W3
5kTBMiXUt0TCH3Jac0iFt5Xa6rpIthirpkOxbcLvgSZMhtwESECep6v0xd2OU1NuxXsFmE7GXuLl
EjT6abroViKdk1YA9mnxPXrbErfbhn7DfktOTgJ19wCvfCm7yaioQX3Z+/Bz0uXFlR7qTrgTSHhh
EUY2llRb6Q8UJt3+BJazZ/f6mUJXA0OL3JZNHlVUpJa7FIszSD3+yzIHotMZhnwnml6kYQrgLi94
xMcCl9hRjH6qoDahNKZbfRUadtj9N+0D47En+eXmWN+wivc8YK52wsuW/Z39plFn3bVOc72ylo7L
nSaWIyXjZ+Sm+jcBWeuSkIydazaNqYyPlBEGrxPukh3gfs4pdVNELJX0a7SGN1a8xxl/x9H/V02M
Zx0sWaodX51cyuMCe+7lGZ2JiJfvSRcHlLJKqLGmnycyD0PrpSCMV8c0ytnMYdOLER225MdhMJcX
g2Fp684JQv6aM2LJKOMYGZC3XYAlxmitwT3W7u2EV3zUCV8COZCxVB9brOQFjdu6TDag6tRotVn7
90ASMKlMwTEIgNywseI00c4Be328KfiWF3XfG6QiNG8bUaNw749aVpPABLx7vL2QdUlohAl883y4
/60RBDK/hFSjmY4OgHm+fdbT+kMjhoBFi1oLJLhA+MtpkFQESkZpCubT7Ctg7NZJrWkMcRakzhGS
vvR+hTvLLrO4uGbj9p+tnYxPbDpAw5h6l1GzQT9odTt/LDMgsRfQv4PbwxsVG9PoMoDxoQi7GYvA
ASaR+hOfIWQ3ObdbhPI/Y3C9tsdvafCsB/KVm0fELeGblXMJSMkOkFlGF6482QqGM42AydBmjHOU
J3+Gfil/vK0rxf9Kf3IHpcMp5TDpTEi/nOY2nEj3ct4mj08I8ETdSgiO/fe0+GlJtDlJwOhTKoo/
qjXWxcV5FSfYyAHKvAqxRq5kxk+XicgIUnIgPCAUYtQysZ/Q+6uHM+HfzXd5EXwGhQxr8A2QLz7o
tKrnA2nhwrYuQuK8sJqk+/ysOiosfRVYi9dBnFPjO8da9oI/IaIsysnTJuDvydPUjySfv8XEmGpM
kvU3gmFYoruS6Du7Ss/z+OoHvRzP115A2EM0mN+zDV6ZT3yABMl6T0AsVlzrXRLA/FoHxPRVpHMK
yOJvAe7dnmDaQhXCjMCAQ6OZXPk28cassZw8TgVV3XOySCFpOwqFw2b6giKAIqzMtCkCzwIjP6kY
+WNPp8+CYylu6oQGjS9aXY4RDkBTa8FNYZX6ST7gL1DE4twfr5E5YIaiCCV8FVoFNqOFlN1hlM4c
HasZmjwAMapxeR3qnNYBBbwA1bOcvnNXi8KCVzU398MD6BINzDXPPVmA4s7/IlxHoNE3KtvQqetE
noJTI/xJX8vice47uD3A1JE86n+bV8wQ6O0WHD5NYiG+YGLyv94KNP1d6L8W97C5kx4G0qE5uEk9
PdHs1Ou5u5Z0JNqFFJylFbrGeEeGdEUcwFBMbNqJTKuQ2AxKWdNxzZT8/ZpRTrhX5T3/qeYvU3mp
zyT1h5pN95+ekEGyuq8Ddu3foBmLi0aqVNIDMhrXDAQS61EflqFbjCvGHECRcZtOOEvzV8yjLbA4
AbV3phnAx5gTQIT3Bffnu43Q8i3QSBKuQfXerxa7xCpQBtAdxS1SmdNyRx7L/hT14zHdIX0X8CSp
T5YyWVbfzwqQRVWDolbOOPpECl10a7EgciulQgYnVcFBakboGG7IIdgDZLck/+aeNkXgu69BZ2Kc
HaTmdalsSj4MftO8yOBLPB6x2sTi5XH5/doW4yYCh5rIctZMEKQtAi6HI4AB3qHn3V9KlpJEcTyq
s4m1Q6GopoP4US9ZAlZYMHDlqRN3lq9uHU+TeuN6KrCWzNy84gdU6JP3jSeYNDVzTuz1EcO1rdbv
Wzw79Uy2w0biZGcKUDUus9BwNsgSOyiJ2ENQf/Mqub8/aJ4yjxhPh/8hu/9ZqTe7JE54sHSJUC6A
CRJz1rNaXTfvPJhp/1SlY5ZmR87VVP/zPc24zNpFkoClFSJTusx6KGeGT+0eqTikt3Rmjzg255A9
CnE30Hox1wgAIr5rtvqetm1L/B8oArl91LhUxyU5Sd8uTBJ1HxEyuEU96UfDJVrm7w9CnJsFPxPf
p0TlHIleVfCP2hL142kevpn0HApaeMOTj2PZSfUgPW9D1gf307cmMJxGVqGYXFr3ixqT2NBJ42oE
e5o4J3ELaFfe/BeaxYz4dH5lzZk0wBudAGWzI0pBVpyBrGio9kt3SbITmzafp1xxqRauRzKJz0LZ
zX9/k/PhA5w9gb7fEDHYLYcrI7fFkVc0qBdbSHGpZGdmHEQjYnqkDPELhy59LZCCXQClN1kWwCBT
cMCAgn/4tbeYBVqUQGpeMT48wSAeDJrdlQtTrRBp52bmTcyy4GZTAKab30gwuggwQJWdoXRRuKTo
XjB1LY4d3YvkYeaqKrI8c8YcZ27jocA1xAfCAawvlXBEGWVxKL6WCy9C80ufPffsaNXfvqyXrUll
PZY37yL/rh9mtDU7DsiQ0kzD7iWzsXgs69H63p7XEhuc3VPZsYJnBnsh3h0UPzXoGTZ5aorLPffy
BwJNFzqwBG5NZDK9zl1mwR1Ezrgms74IlFzEejH8Z0pXy8eYisRJpaVf+3nQmVd5KdIGBMSwZOq5
RY0jI7cXvYsUPpcP6u4qKqjj9r83UmNqNkjX+/Ax+SChdQThsNtMKxi4scrXv16nrD8gLDL5MxFz
FW5bye+pqO0vpuetEe6r7HWkcbSMT31iNTOhDZK+zhrfUXP1Rr/n1RCJssGsIsje1azd2rlsZ8Fv
Qty+UGeBh9zop6Vwp0Iu+o1AAOrfwOfdKbZM0ApWPPtEkmTnkHf25a4Whzuj68y9UXB+gLA0mBla
+oqxM+KO8scVjiQMql3ZN3z85ZDnvZreldcoY8+3fIg4jxHn303GZLyCvaoyP4v1IdXa1q+KVTZe
PnucNgS3io4eqPgria8kJTNkIx0fcJCvcjXUD6vFjiVF4Bor4ptLSNvWUD8XH+XRx0g2gsYObT3a
t9ILSB3FryBvKi60/1SnPatwTSaJqEeUddBbxPJRQlC7jmaIgY0+Cjm8hZ39YDfqjNFFygm2kYBS
JIDxvn+9ggGNq9L/ppjTUtjyQRyQo4XRene4irmzfmzYNAGIgIff8nk8zGveaHPzzx3SPpLwMkiO
krvDfPlb+0NCnbLEQbVFMsfmvDTpNDEE1dZxmNwMH0FpeaRRVD2EVwi+X8nmWVsTSHjlMqFut8ne
UgSSxESMMZOlJGVwbDDECTIkswx3b0Q7r3rQcbdxraBKuKw4/DvJWMJi4YAKOSSVSzBepOwhGt5B
n3vf1zZNlhdWUeHGWBdKZ0SpNyAaictAxGusFx42wLPL1dgehVxZyORjjLUKG/9LVBtMt7xvDYsP
rZN6WPuwxjcVz0uTOsjkN+sNzccLlpYwuAdJOT/SeZNOUxqbfnWkm2FZ3Ldcltr+OjVApHzChxmP
3G39hvr81UihKLZTSqJGlLhiYcmMCfS0vwk7GR85UTF935N9/oKsq1ifW3eiFPTnzxiU2HFatQZ6
EW1X4hp3YkRvUaKQvLXG7QbuHdnrs6g7Pe1uo6IqTTZTq5wy2leE+KR7+yl8VPCy+sbfXcKBYK4p
4gudLQN7BDNJLJw0fJt8R21cZEyra4SvY+aTfA7VBwHfERuoEJ9Qq+KMHN1AuDZc4MPr9kb8Hefp
PWwRnJ/ro5/Zr615b67oOC36M7tsjOTfZZVma9GcR0LlrNdS8Hl6zur8XkEs2/IW8i0XCEqd0z/h
cXsjJMyJ33zfbRFALYzho4/gLblPLbKaWWr94svmE520aKZxfNBuTF6kAXoLboFxXA8ywK1lZJI7
TiR9dF+q72SImiAO4Yfld+QGXQC+ksGJjDZlwntOeKkzCz2MgRksLDModuJXiRgdxHQ0EZkyUpq6
SP8oDguoUfbAw7EM2fMgGRuZ3k2EcL0mO0ptF9dtK1vUz4jJnuIyYVq9wVRZ0h12lzGx9A0fPash
biJQTuMyBT5ZZak2FkkAD3iT03eRKOunBP5nLJETle2Nqa5OA7bBif93SBBxRawr5agWo+vYsC8m
ALqoiTR1QiutlfxRe8rYWUICle+T9t+VpZcW83grdfRChkjWjefGDHq98anLl1aSkMgqroSKNvOw
94yVOOxOEVZuQEKDO8ZwWEeLMlHCA72JFwAnoW3hTzc/WdOSrv8/h1L9Dx6PSKscq8hlYRAap2/n
irBivNzpdpisSECcNoCu4I0joz8V0aszepfYh8ypYv44ooyLBPlXGofuP/oiG4kYy9UwGLUi60BI
p3+a72DqR9hJDF9t2qFC3mnFXeK9slqk6ILCNQKpu0lmmcWsZpr11EDkRMf4eGE3os0jxHFYvGdu
wOYZVtShpCGvkFdvRfWVTMsJVX8KrfW/qrRoC4FfuS6q8k7w2Gbx0aEdB6NPEEcoZk0NrHZpxZkK
eLGf67t92qLhFYlR4EXRaO0NZa3oeff8WehDtZmuhkWDIK+poGWlML+/ImIJaz/qXPlkA5SOdyBc
Omfs2vPqrJnQ8HICaV/72N8qzNNqI4I6G108k4QgURT8ZA+bJiAm7fcRGqdz6Z/lQfyAvp2IYVgi
HeMoTF5NyvgQBZP+IwOgAEsIVOR+k/jxyFsTogrnfnGUclMhpC1lHvUgj9icEZgc/3yCkLMyW3vA
Pwmp//WJTXVzCjqDxxiSgh4pAKMWnXFodlwaomBrwb+psU41Vj7i7uU9C9d8GoW1rFDuKbDg7PmE
Ig1tIaD7rEPb6unqGz9eh5yxKjG6chOFxfwfHZDeyL/GNgNmo6F33pnqCBkiJ/DBVPxr9nmrtOv7
e8ha439OHGtLPUfNfwlf2+TlEHOdHROitvR6f4rSN2fKY741RSG/8gASbUh3EwVtuYbCmxtbob3K
Rkk3acYU3CK4Jv0AC+HDNoqzY1qAEAPtTRpBKlgW7tzRv0fvg9cg+XAvdDV1oxHp/6faXOs281kl
ZnG4zS+NMRDhp2xILHKAOJK+xDuAVTwqh8gUHj/4yPNodJEsVbDkpe7iIzIEdj4rtU57GxrBsS4j
1kbQjdMkUeRXhE4UdoxCNPzjsl3ZZLdwn5VvMnq2XW7k3rBmkh/HWK2S0GZFJgIIT9uJPODpH2qe
aw3pTi8gDyYv+FGNKCSkZDmp2MqE6iRJhOigIHdq2CB1LN7DZ9UW7W5GKPv2VXTVkJ50vP32wXqb
BupRhkgD3E7DmMqnv23NowKwkKuoDv+GIVBKvWbrLtAy7ZPpOl5K8QZOviSiV+mIudAKENwyKCKL
XN8YzwIwYjZ5SbAH/fJPdrtS/sfqAQ+ZcH/flrwx+eGzMWWmJYDppvqR01ixwmcE3xwzFmaROM99
lyxBX3c5pBC0pbUJLKW5qtszC4mewsCHwi9YC72gX2+AfTAiv2G9TaPPOmkB1q6QvPycwMZ2AOIS
YLp+woB21ADTBbvVA4zyeS0kdWKuvh8PjDb3m8b1jQYuhF4XMtuAj+3uWx6RAbiWUNM4KNlVum8R
ipjm4z0V0vx+t8u/yDUuAiisa5QNFLzvOAPS9MuD0wzIMgPBzReZOneMR8ATMo1NhK9kcP/nMB4A
iXKJ/efWz8XvGfirxaxWBVoxJ5lnSvLhK87JG4/YcaUINi7/4jkUOoykXLsvEIggmUaDR8woK8qx
Q0qgweBetDLZOdAkzEmBmBF2wshE6ui1FgWNzrwu7F19VDUmWi9fQKGqq+IHsmpf6O+xsIDjF3QE
WHvZYPtnXrH4S0oHskKsnr2KiJKecEY75h4wFCUWe41Agu2o1D0flHAFTddn3GUlofIFBcKgC/Sg
3kqcc+b9EqdaupQcS6UmUJFUGn1Ufi/7uKe6oXy/CX8ZpVwZiJHjMTrQhKXdruhYH2zxVPGJlP6J
wm4vrN+9gEy8OoGVGqddTIH6vu+jvOCdMbT/wGXXn3tSdJlOxQLOxgsd+bgXm8n5jD3xtkck6ikG
I7FayWQmTw8zMTvnz4fLF+jNFV0nkNnB0HVRDNgtFYYKFvDMBYBKtXEJCPUwt5QQnQVtTuecL2Xs
z9lZfyyuRn4d08fmis5Tx+Tw+Q91wt5IdI4CBpBFS9c73/CKGNmL24LJF4PnO//SqsT1fIJsz2ai
eMTKOAHiVwxMLGBf7fRqAyPiGL3/sgK/LaanIulmvXlSVtWfmbPquLs3NRHcgnjdbwxdFAl54Nr1
yHZu4H/MNO1i8/HoiNj9sH7zgeTWlQJr+FgJpxETbaStb0xUCE3G+iStwB/DAaWVK5j6NGk4AP4h
mPRlI8vp3XMteMmTUDuC/dp6RvMA62FeZUxCrFCz4m+tP4lYbRiD+VuO+GxxdLLilTqYj70jQof3
4WrZtb6ubuR4n38EJFsB4lr72gnduzrZXx9O1/+pNuPZSnQ6b3W6fgLpsO9vJkRQKet3Vwh33eWi
NDd5tecNA5hC9LV30+Udv6lIxEbrVpX/5eJuL3DzWA9pgyscORQnZSY42d/vseeHWRjMf1sKeuCA
9xtCnUn7w2UR6EbdZLaP3IkKh3aZVLXI+jpj4cFsZJ7gohL9mibuBBUQ8RB1AQfEosgFayeOgxqy
2DggUzv3SI1359iriqZwGb3C1SSO4Fk9fMgVKEeHvmkY5S32DSuTMkrCImeeahUTsZXKP2nY++nR
yl9nKq95l6veiXLBprAOU6agyxiZZWo7bejQSLWT+GGrvfTM9oEr6InuIbqANkSyYUwdDJrZdtl+
bXXsOYJfCemT7J8l9aWIlmXJSW5biY4B5j/L6pbV+D7k49FPFhP59Qkp/7WaQP6AHvxSd06dVjmg
OwIWRH0QUHu266ZwFTp7AoqfToAazyXKHFQtwoOG4wQHU+sEtNbFxS3Shpdt4pIxm6fUu1sweGJA
JR+xuft2zW0RScpqUPz325yaqx1OWXCFGXsR9QkjZdhJX8mfK5LGEaSbFHx6HBCqwYD6Ixr2Ket/
wnFmeQc/8Pf/Z2s1Ti/RihE/pxx4SvEST3c8KLdQ9WYZ9qVMTycpJnNWFQ5VmlvvR7k0iDYd/gtE
KnWjVHH2eOW2JfpSYwFVSuz4KuDx84qOU3NuN2t8jZ2ZlZOJqu8vbSXBeaJ+uRGlk/re3rIZgtJz
3WQNj+hm4TVKaFh9IMzCTTTf4L+K3XSjBGpFshGP70qQfUX9JoUSS/LF/Qzcl+3CmaLVH6guZwZ4
/pArWAG1HSxUa/XPKcbkU5SMLgBj5LMFjbDkldtZ96znqtyxkZZ/G9hu5wNM6mXKR0HPuY14rSlx
A90bn0w8XuFOoqtoV/YCJtoU3eNcSM2Tr6AgPgBnFnZfl1WwN/1reYDYrksuigjrDoWJ/3U/bl3Z
ji8NGsUBelbvCTW03oaVc2O138+JHBRbOEZEzhkjGRUenYRFpErQ3SuCePOB1DwHDrJgaBY7SbER
/vbVrZnDL1hv4yff/gANNsNzg4Eq49lvXKW61OIRt0t5hE78YQwplDo5Q1XEuC+vvK+CWFvWj84A
uByEMPzC7j4GA4oHysXHFJlpLU81kHJ0yr0zlRLxSG1oDbU76ayO6TWfYJwiYtMIsYi2O7OXW/DY
2ATeooZLPoudtmfMgCS9jO+GUW+8HiQeHNbM/B614yUPjIe8KlTW421uZML1ELrk3UxA249vekPb
YUeahwH5jQAmMBIlzk6rYp8lZ3b5Hy9wWn284lCChQE4KZNwNEUVDcUeYwu0nsVmVrE06lTVuW7G
vRI+OPJnYhacSmxU6tK4NPOw0N8dqmBT+nL57Iixuh9Qfw9DXdPFMd+XlDJiJVxi2dsEqmTOvdB2
Z5PcOajXO0zF59BxF25M9oRjCwF8xgUD8mX8lzCdTptBo/OhUiHtk40jgKuznvMmQepwmtDRampi
GVSGuiUMKTX6/6Ssb+fwKs2NqY/2fqzwlM3ycoMsfxei+pAg7iJ2c2EEQEDMIp56QhUkjK1aygJF
neRN5A5nQOlYslgjUhYdvwvZX1zUaY0I/yJbw6z1wD/Zc8msesKDqrTC1GVyBFAz3Jo16zsacgwz
uUTI1/oS26b9ok+XLrOIkjk47naG7UW/FBC0Mw91JAp4UnHnEKiL/tAWCiA/cj3HJkODjq1H45v0
HfJVA6JuEOz4dgi0VRxUq21hdD5Wc9ZN1j6HGwQHf4oYzXzrvSO/miQmfhgT9DspQsXu3axTf5GE
DqEbkJIfZN8ehXHX3TieQZWpfaGXH95QquiePDJFXLGtp9MurwIMhA0rj1QRhm9yroBuJQdOzpIu
0OERf3mE6l1Ib8VVi5E/mBaoNbzLoYgJOvGkZ+yR4PnFRTXH96JEU/aZpCmhdAGALDhCb4VJdFA4
DUAAbtnttDnqUp7eUBGjFJ+Fl4rTJVlW0oyEVLowQSPngIigyxgeHqN8ShVgbDNxl21ofWtBL3sy
eoEuiTvQEZ13yrgmZlubIgO8Vg06dco/H90GJaeEChZlM9RorLaIYO7VGNWfiCJJFD9bdg3cjlWn
wCJNbtPUAGflFJBzBb1ruyRL4lkOspVUb7EZ5DMuv/0/KNTPbq1Cci5nsTjw0+g9djdnntClSZgJ
aw6PsXVqEhz3fTttrMGQpLiGeKD7fJo8hoAjEP39w9ogrSSNou2MzC+TZsu6aPpdQRW3lM1s7GD4
XrCGb+7QvwGmLrFV0CGPggmbErTRLerD3HEvGRy/uo0pQdPin1nvlvr4c4sWQROH3kQBX6E4WxOZ
asU6YnFc+qOXx3ofwlXHVgotX7UEcJjWMt/RYfzQ7zMMod56HF1SPaDR5I1uHZMkb8l99xKMJdaH
lAPPI6ZoQ4hyNHC7Rpx3RbYggXhdpcj74voZ+jnoSK/L84V8bLcUfnMX3qfNqaAYKmfdp8wudj5b
+iDxHg1PYlq7Erwf/zg8wH79JUr4wrQtLAOFiji6W3C054RwyjNm85vI6nFcftu0koRToqH7p+nk
OHzc+Vx205u+h9oauuF/XzXnuRqqDDewF5hPvFS7bm5cH0TAys11eqgY4SmeiTE8JJ2+pLph61W2
4ZKpI4sEj1+dHfb54fh/kbYugw/8CH8/x+k0LI62XrycVp/Xg1NhzVlJon7l2fUihPO3IWZmjey5
qqRYOmPFBNQiHMCrT4WR40balrpu/S/BKZCdrwzL6/TJVBZkRh3UjAvadmF62Fi4RzRdPnIpEgeA
d/s9WJJQpwqtfpI7KEKfz6L0Ae26mBuKVhV4ZcVvw4zlsLnLbGTHVeg35yZYHwP9+VVRZPfx8knw
bhfWM4/q9MWtGnAAy/wT91q45GBFKF4okkAvg+NxAoiF4JF/gcBktS5YhSrpEJPYts/rXGGrPv4d
HtUKcU6qm1THkyJ400QhO+Mo2rqVN/0RbuXX/dooqnDiizWheHNZvrpe9HSK1Tlhvzq4Ifd+dKgy
oLGfB1GZPXgR0Vjg4oKxMlhwuFLXCOVVSO8SkgvlFdjnoS9IhKqNejxZhAqKrACR4u9GXSFV8Tj1
hsb0JnOsTPA53/TzaVoIEsU9Nvelfc6GhRWbDf+9kQEIr89qg52P8JMXxySFgOcgrWb5h+yvriyq
PTut5euhQuHeEBCmMWY21kSu5+0WLBkybE3ZJajIId2f55hoRB2TybzEsQjNqNLvvsVI7at5X9NG
aISzbRrHtchyrNzvGAb4Vo0HMh+Jh1+JckAKuy22+IOgWikdWho7hH+SEzmZE6GH+TTiOZfSUhUv
Kb1IKOBi4ScaN9NMrAmLIG7X0/nUitUsFJFLnbb0U++8ZArZpJFGznkbVDlkFiraIzypANKlXheN
KYewFHBc/rrPEx3qY/OQDVHIJPYZbwMSZTHtwZAC9X9a1t4G+CW4G5SXNwslCA5mcwiMijlcynN+
8Nqd9Um3Fh7IICxsRXStV0Ng8uxBXdn7wda12Rh7LAGUmCoseyi2tZgBaXAVcKLETIxWW6PC5/WV
Cl7gg5qZABfwX2apS/bVeXwyqAhX1WEz1isk/e1Yo0OBrp/foVDAtz4thLV5rwdpIGU+U6FM+YHM
50w0a/hJn0fQ/BHAJ32J7TShHtfJ1nJl9lIFziIW3vNEA4XGSrBlI8eaSMEXoNrBMOUGq7rUjzgN
goRXJQvBSgmWBkHMYx22gixkK7H4X+7Zi0aNA7Jg93ro5XDUn4pzU5wohVEJ+XIakJhxvrTAFZwe
jRK5kDXW0mHWRpsMclyiFawXa7kqixfkFrqtMrsqgB2RdJy10f29dLv6x8enL/Zcdfw7HkyIX4gK
q3iu17TUjWOPKwwuaXOh7Cz5R/IvaPbPRJX/k4Rs0X4WLdycMzUFPMuFTb0hYeZxmcg0PqAcIXIP
BH1HM6qdCKIJfskgCPOcBuyfuzC30fW5AOAo6+gWsvveMlSDVcnhCdHr0R/pz5DLP5ojVNwW8YkJ
1Qa+r/N6VISAFvjhJIvU5caA1xYnA3IiIR7g520t96xam8y8kbtTBJCEDn27nEtp1lWubevBDKJi
zqyb5zqgAHRj3w+VES8hqtNi84RlKzeJWYcdNgbSJ+YdgPfZ+8LcP1iJ5JcbzUbp+fV/Nl8+5ZwF
Q7wMyZ+mQrw32cjJLjbiMIMMR7l08cHWReYtmTD36m8Dg8WW9HP5tFTfjmNVc5gfKeLp7x7R3NCC
4xcNGJNTQZ+X9Wt5kWj1ogUCYoWvLzAmqaZGqVdEFR6YrjYT3LHp+ZyapYOc4X4i/JH8OzeiWIpP
fS2bdzKkb+24HPbKgQSjUV8V98cIiv85NFhvR9AOwT9F52eyIbLz7Dr7JjwOFvnpasbWns7PtSpo
S99g09bjpCW8AYEIumlg711o0gZoFULm2+WvqdkRBsTImG9UFBQE56EvvWR1M0jbeebqyHzSPjEd
f2hBcldAljWZwirKD8aJ1nWfD+9V0Uf0KNxdQuBfnBIAGdustOXpGxDPcwUIfChtEoD+NQRsVhox
Qxxf630Wm6pL3HYiFFUn9JtflEPCTWmqmeK/TTDNpvreY5wxZTr755ALWDwgAuFmcmzluoIVicGr
5h/oW4sxpXa+htiOYqRwweSk205aBNCMSCWCCgnb/wfegPRn/5Ru0n6tVrm3NYInhTTpn9OlOshU
NP2DXKxXGrOFO+Uk8WYcTnyb+KOdq4vd2ByakLWMHPgwo/wl/TaBxY6F2y9Y4jbMrJzq4JyGBpLm
yXnQIJ1NqrU1i0W76EteRCBhRm6TQ7odwatVMN4B8Q7hhW+95U7/j+MBrHyDxv+evLfGeZnjPx1v
gbO/6fwhI8IquQnYvzHx7srjkNyGzmIl86/DL/AaLZswpQc4rj7Xoxx9Qq8E7qazco9dtKjzquk6
eaNPUu27HIkBmO6PmK109t+vQLbJU36OwJ1Yrk6UosdbwU9FlnCVgzrSxeCGhCNA/QA2R0C5Ddei
dZBclhwYkdJHcREQhYxPsVOUHtpzgqvo0Znh+nT96SnyYxHMdy89NmWmq1R8Y7vgC0tn1/nh3gYg
joss9qGSo7DBExTMWOwmNB9ZgXtOzl5hjYt4CaASRNvmZfTPEgXXF1Isd6beblZ3CROSEZ6x7mk0
/DX/ATSW426hHvSjHKdMCeCiSvcIcEV37m7/NTvZXIOnG4c+QkB+2AqDGhEo5q73pGswYggNBAmV
X/MZsm9znlnAdpD1wk4S24t0cUKHNrx82dCSke7cpkL58v85kXQJjmWyw6g7gXV6+Qq8jx8BxCz0
DKE2VqAbRZDhH5/QelE8WQw9Ewvvnq5vU80dXDP/jt1mz6I67AMbpRjRIfkApIJR2jV+Vo9a57/C
2QuzeEQSepmtet91ocbSlz6LCO9YID80v+s52rdI4tbTYDA9j2X1L+1abgN46ePFi3U82FRiDLfS
yfjvasYA1uYpW/geeIvNTTO3CnTrxICXTNINurq99ZKDe7dffSKrZSUSykeepq74/80PCHe+XiZj
fN/lAEQj2ElTdHCAiC70q0ZeprRapK+oAtXgSV5p/yfgLPXCcsIksyuqP4BoDYA5p+Eqf8l2SaM0
v3cAzlTCTMigq6sJKD87XEMt7/TkURgto0bvS+dMzgLYjzCbuzQXtQjRbUmKqkPm4sWGFq8svbnE
Efb2J1bcHe1UdthYIedTQd1tpNT10RwvlCtZ/igslwiFpI267yuNmx9b6+2VR7luM4K0kvMXe2H6
iRGH970br0qDxktHHWwDJf/6azXAFYj9V8g4zHx3FT/QyD5JEG4xmial+N4aOL+aKmxo7X8qM5uq
Z39wgmeooSdSOAbDyjO5xB4QNvOUdZaRAyyLdYiTn18Vgff6oDbgh1NB51jcv3AUyEGoteGz/1q3
4V+CFccKG2ohqMidv665LYskq9J3pAv0QpnSgx0at/d6Z3tpwbaP4qB0dIw+7/tU7w1uX20OjaCi
atGtCmYzssI03OZniKHUtW9E1s/tnrrC/+tnBOeIs+6T3Vycrwt/OpCaIAe3fJPh+wtF4IfsLPCi
y3XkthEYA3miPZHaETRL4VyGZI4tHrmqWmD+vbUIYIwujvm9Xsung176cFP+uVptJzLAPfhktezW
fWb9MGZBwpT1kUc+BoFySr52E7TlF7tqywX0ID+/j29sgckxCNtxC05EHEkGYs0s++DsfrFxqXgO
a6jHayAqjcTbpncrLdcm3rGqlTsdsjzJSkBJ304332t2ImMQIP8VQvCH0fa+Gok54Alx3PrbThoo
hP2Sr49RCPx9NBrxrq9EleMZcL36XQbarD4Dql/qIerJTBgIqhnEoI6or7kr/UtyGVW+VCNXBxt4
JEO1Y/2tk41KhvpUIsxHH80wTyeY+YdM7bS/yPXYnrhxaZ2N3p+b8VPtRqZtFJdHrM0NS8fMUCDT
p8aw4bGQggaqUZ0A7ZbC6wl4VFBmXhJgk1GwFLXTLdBgvcSQmQJSu6BLS0gy3r2Q0S0FZe0x200C
8ZPn7xDNKMKi10IVjEewd7SsZLVhK6EIriK69htUOUVxDoUd1xzwOK7FaG9k0Wgoemw5esiTPPr6
3mYX9zqjSSOdEGQy/mVbwgQ8FRReb5YmrSRR9KJtgrx22iktXmHpw2cKYRQaqN/RQxNF4keB1EfX
2H7Z4IFhyj6iPgss3LNai6H7sYlYeh3XtiFSVsKIP0tcLPXZgElvhPUvc5GrF8d6Mw6p0rwTEx5+
hRdn4sQdYwFvwNqJrOijr6faVfpitrzQDxI7iFr7SOjLw0uK8FPG/gxysALhAyrEG8GIpnS/vYGF
fjdfzMk7Xx0OW1l/IfTHST0M6BpmOyuhMthXou04b0xzmde9/7Raa1V4TSFhGwXgMBLoIm16Aaev
tOOIvwicy0i1ptgsqY7qMqeq/TH+yDYk7fTc56Z2u9gaf0YP0ClXXNC9heTn29uJkffMaIe5x0Ee
56N3zj4v9pmPH8jU1k/qHFAoGWNkn7rGt+97THeSEjNZbxDlCpckmDr0lffXOIxPuduNXIuviyvq
ik/QASVkiYnxTF8nkRcuguT4IcOSyXnHsGaNHlL0W+lfevWCEF6MFj0B5rqR1thPOhFS5ZChDEgp
ocV9QsSd1IgWc7Mg+iC4pKJRtXy2oXaL2ID4M483RYZaQX4UFU+6TlGDptUyEd9ueloMKXjbNOOn
KZk6RvX5ewiAS0/YLbrByEeIOe4zlf+9xWnbl8+cg3MNVntUyg1om858qyGGEi/et/jkZvmA83Ar
cdSf9qLueNzRBs1BkT9tK7/SMBza/D/H9RJat/ZvvhRbTJ5ZtSKT+XDuaHr9aXREMQgB2KAc99RK
N7tpUVMOQIFZLIryu3zuzFP+L9fbuvHNY96QFRVZju6pbgA4KosA0fvZOCLVVhamQVE7hcVFqK2I
k9VuzM4B7OHbCim9xDtBYwer1jx8vI+D7XyUB5AL4CRXb9Iz6CjGDpK1D4mLHZe7m76Ahe11uGGa
vzHSEZq6pcZICYD6fdvaGEKix/yakDYRzkpuVoBUI2TLL77HQrjeSZXYBd5Y5INFJGk5lHHq5MWf
AnuF9571yxXmEhZhygqe7Oj+w26tEgD/d6fA8j6mAbLq4FmMUPdd6DvX2KI9+J9DcGBAd95tc9+H
1L/dSpnWwFpBFRq+IyiCNprEfPNQ6P2/AIHYTyKsOpaEkQHTol3CWoUyD8hWM+Agi9EgA6ANiT8B
0XUJJ8Tezrkjw6oRMAhOI8iRSKvBO9oVqOv6ET6ZJ7hqp4gfSv7keU4yWXkbobVvGDZyl7Zpq+t8
GCk5zu/dp+ZCeNN9bURAz2BIN2e6YwfGLMwPAmwqSeKtHrGCqkhL2A7x2b1aKfLyGDKeTMxIfFhG
GePfBhqfNy0Vjyq4nSPUzJD44/Mb/Y22Aq/z8RaPZCFpLdIGED/Y+K/I31pkLNwlXMeuE0z3lTRG
W/XqVfB9XeZ9VWWTSqq+Zhoci+BZTQSQmUKFMJmzirf6y+ePbDcJT0Zo6XS52sK4xV0WQYG15rW0
5EJw7fWwWlJ13M8PpZCrZtYPZPMIeVSkrMDXEDberhngeHdswkzsZvVl2sLozfJe83LjVtSlqEck
WKDzDKWoLP3/xc5YZKeXJY2le5ayZgbVsmL+5m2NMaso1IDmhqoAgbC2tJJCq9ZgKAXrAQOvvdv9
VKUFubgcVc7L12mI3fHLepCU6Rplv7gzzOZh8rm2v2DskUxcChheUpFX8c0VXoKGLJG6wBFWdDHo
HWqBGXGITfMlIfWldx7yAIUVFzXkzeAQPMXAOrgf9JzZiFwvpSuyMj4dFgvCD4ltAKi7B8zOzpq7
XN7JTTPgUFLGJcwnB/Xy19+CCaZ2CLzapgYkQRv7ew9YCfOZulpjMUYRPxiQ/G73RNDtup7srPXA
1V/cwtYoINbYFRGWAc/8eCu3t6kT2I31rabTLaxOrF+AJ3Qa9fdVjiE1SwStYebvbXp56cVoGpEc
/2d1p2dMnU6UEfSoy4s9Nx9ZHY17nIZsgZ4lwWbsHn3dSGybKKNqpRsgeb25xL/kis+8FVQGno5a
axv735crm/h40/us44cVPYeobkKasoIL7R2jID93hPhF0Pa5QPRKwOFtiS9nQ3ZtCzY5uw2CA6jV
z7nOQyeDpZD0uU3hTlf/Lv/M80dTmYtxrl+4XwtszUpp9swf2URQ872BgBEWU5qXJuhLF5qiJbe/
qp9UvAeXb3XI/MlT+/pY9LMAkQ3K6cdEFKLjKmnWbaIhsro/KlRs8AAtJuhlE4+C8seYnNXIWflF
L+fk4pXF4BnnTBlUsDs9DmGZwW2qBqO0OxCTKJd1rP9IaplClBCz4B1rVBxvOwcEq39szs+iXlu4
Ry3xQAlkBx/e5kkXFxM7yFXg8GRmiIO5tZtxaqltA44sPdPV/4rcxbifnXNPLyBs6PjRQgdIP+/I
i+YGUH8ZFejHO6U628+8NGAXRXNPc7OF5JT/M0ddniRLHRrHcSuzzoQv9n4lsHjuD2FBqzBkVtf0
ycMGnapD3uLN84w21E+Niaama+bwRLmFfXi33GuEFeaZLQrtdQ7xcKmnjxa1dZV1alRLr0eQRM62
BTy+hSH/4rJTIJOykkWQOfsG/8FRi9+X4pBNtXwjail8T+vIw4+RserudvgIyBwtnSDaro3sEqic
nKfS62yjN5Jp+cFm0Nlwy5cHs+qFBn4zBk6D0hObK8QzLjstSCQyugUW6SIGKNTTmbQt1Z4tDdHU
8e3TZpSwcSfnE4h9U20HZJzGMd8RcXISnkK2FaBWNU32q8v/Q0KR+u8UeRLchezUnuG+okM8B4el
HczxIU3U29n79PH5SWajReVmpeQS06jyWdNOrkYuqaSVrjZd4BoiMPUAeKh2xOvA2Xof9N8LarCS
aSW+XYU1RAxdT+pqKa+yjKwpLgEAwTjDs0iQbWD1xJ4Bc15TcpRMaW3GqXGyDF9GzQScKGkIWCXK
/1MMUk1izZXJtSouxLrFat3uMaOEv8RkgIVhPRAlrMpQ+WI4S4kuLWTHH2HdVH2CDusdPbaYXSU7
VKraa931j+sPnCXv+nwHqYd7vkVqUV8NOQyEa9KGtiMhCbIp05dAgXHRwEuYjJ/vT7ph8jNzVBDd
t14cDWAX8bSJBbmZGmFDHlUwe2xl1Ui+uBhJKIZnEi3D00aBTvrkwkw5+KzvqhdTt40CH8O6qKdp
+tgDe08s5GwDOOji12seru9mQdgP4NgGURdRSZNtwjw8XkS5acn0jfBv3GVHSC9WcJ51o9sWabTf
VksyqSeYA4Vn/ObbydPcEA34Ie54KuoW14i00L1s4GZvmTDMlK1Mf8FQ35jSPow1yCcAJ3M2Q3NV
hMula+dSJs5yps0IUpWiMtb35oLiNZ4Y6ScSw0BClb4ryLWfLyksBurbWZN+AGElCGd3z4nQA3O1
hbkDtCj0R+SigjHv5K7gEBCn3qxAFcFknfstR6cUSW4mQcAAFfNhmWRV+BWahJ0hSGT9OoKNbu+j
9PZ3Mx9+0Wb9SLEc/Rl5jku4Eo+L1Shafg0mYUOnvwZQsBSny7pTIhqdCqTiNxLFiEAfHTm45kZz
jRrxWU5qPWcudwvcWFLlwFmZa2+nTpZ7hvqB2JJHk+jSli5ZhyTNomN3X/vmVYcyU/qI8TmhMvM1
ijyHBWZXypPMwUudRSUeMhbeb4XrAaqsNK1GlBjt8WIoOoC9U/5rYb00Qog2B8stkz7aGJEc/bzg
wpwr2SSbClaxw81CxCcMUQASzUDAhCEU0w7/uo1pE/EOfSiiAPfhMHNWGC9rXX9Yf/kH4FhVVpHv
TXQ+/2pk/TE7/0eEIFEib1h1ceofgMutBqaBvmA9dK2bZJzS+0vG2YijBg7Uv49TbKNV5h8FQC/h
EbQvCaERVwbfAv397X3T8AB80GmPRieXrfUGHd2hrfUV+eyEcJ7zHt04luXviw317frQA5tSrmiG
fT6qpksCi0WaWgfrhTmIEiIh7un3Y5bfniijJe/XEq7bvjn6DEUKxf/4QuN5kJE/8mw/Y5mBH4vh
ZjO7VdR0Dgq1XqQ4gTd1wF2gqlp9naPbKtDJv9YM16xJgX9ARzwYviQxko3ltf8I9sNc3ht8G/XX
HNTm2IFRdjMy/WAWqzhHf8lfcFGOwygbVsVAqcHvSF2f619c+Cy2hWKe82vv5GSDW/RYN0y6r5zJ
GpvSFOaqBPzJIbZAbpfcjfTldIAsk27fyy1cs47AgjbQAzb+1yC9YZWbtUnF9SKaMhrzQPwYVOUw
Studjv4u7+ukIwv1IeKh8vWbGOkMBPgZ5N59TknQB4WOgRkzRC8QdW9Nr1tSXn8cwtLm/7MeI+s0
/KRLIV5nIIoW4BGX8ZIRj5Op/s+nURWh01MGOK1eDiZWxVXuaL2X12AijlXsjbNpdyCedF0AFfw/
4u2QcY7o4j3L7R+yM2wjXIjDfNSJ05zwxxj/aBZVYNlp4ZO5D6a+Yr7skwE8BF40raXQvH0UL+9V
7ICJF4zWgoVpQO2HemvAYcj9nzKn7ZS0OTCofCeP6fHgxVOFumyJ+pavjR+qN7dI3bzzDpqVc5+t
IPbrn3eQLDIj58YIoXGDbwjgbc8sXoJG6ZKAD/zT5ctwc1hT9hi546sEEMtCvBTeF3vk6IEYpVR7
yU3sqZlqQWL/KgcSCU3zP5COcWIkhlHr2U2ShNEgR+LDpL0fOzwIvxe8D8ZPDLGLzrKP0C06zyig
hTiTS3SJuebM2iHXudkf4FSXucCf1XmTaUqjtMuj/L2XWad4gDOXDqKEueYbjcocvAnA1SMRe1kJ
2eGXZ2pJE0RoBxVf8ZK3y1rBGiPM/qHsufLl3OSZ84H9x4a95UwikMlmLUo6pNaMAZUaaCa5nPW7
dSa1bQPtlmMdtiOuClR1VFYd/ltp61OiHW4dUh7ikgf7zRozpyWacLPcnGFL/5ZHhx++9t0dOZNP
cIKiuFTjO36xDQ2PAXr2iCbBBptpDSxXkA9y7NXzfeCapcORHKYAzYZ+1IwDusYHe4FQRnLw25o2
LvUWHP/387p1xdqhq/X4CnOlkD83QYX/1mflXkpgIYrWK/W83UoZNM6QPULkCHjkQQvlxdI0fR1h
zntwFdzvv+mVkSJJ2TalOMvTpJwQlt4zhN4gJXYlVkcj0/blTUFTn3TiyqFaCt1m06c6L++iCwjb
AevLop9cLWm9+HvUs6AdYGT+HVXdT1zliKuncyuYaHJs5xXxFPE+579uykXF779VA6mUa4JqUDv7
PXpy1a/uQ87fFpEJP+K/1cY1a6h0O43CZ3dwjI1qxwiZFxeSpeGbtSDIJ91De795KnTLokeNWr5I
eS80cvFR0YOTKlUG4DWVu8KQf2NmuO3y2ih4dS1/XxZAqBjETY5MqYBx8/0AAANUVXbK7UzDwiM+
BpkMz1FkaWPFaxMKLF8xCfBZEaUZNIMWkxLyAqxxBOst/MUZQQYVnfg5IPmMdZgIeM/L1x8WCQ43
ECrne2YR9jf/WY6rkbfKdmSLetQy1QDcniiixCgvOmCGSQ9IPvVsHBV4jTI/qwqkobxmiDbFggo8
VQrrYs4Qh6zPmB4GJLuZfkO5T3a+rWkj9Md8FqB/I/6Z+OrKX9+eWYcvm+raokgLIeDedXBr/sAp
oZuRvwx/lZjhtK+oahcGY/yelJtCaNU4RdWlWk/f6KPwNkF/wYduNhiDIneQj8D68YJZYvPNNN/a
sUhPwB3tovrunrmJ75o4PprQospkVbFojfICDIdFe5/bjKqbExgjNb343IvmQwhgAAbHpRMdBFuo
JV1XSHBRpE55K2p/JZJ3Dlwv+PEK8Tc0L4FSgZtLW3qvADG80e0whmddR9fh0Bfb/PR1AHuaFCZG
VZdpGi3ITV+U7CSK/eSCsT6EtGD7Zoaa9T8ImsQ+Gj4sU5xNT64i/hiEwY1C5E8Ximng7ZNaU2yD
/ojjsEILyTNaLPz9L+PcCdITolk9ESQG6OPy7uVl+7KYYji11c2beCPHGjlCf29qKOHu07GO8rbX
zg5dpjuxJ5dYTErZnaKqyuYiJCyUrVxRPwvG56lHscIe72Xrtmjtib41miYzdS3sMzmDrJqJ9uSk
iKquVQxTzSjs4CPbYAAsvTfNlCdV6aSr5NMbDYZMkYRHsJsBEYXIo16V+ZI4ljFts7y7DvcKlpqK
9tnTdsqRe8+8MtlNxObvCLnYQR6mm58zoN13Uvqbc9CMT0/uID9y9NV5DjAIrY55S4VvDemvxXbx
NucDdg1tE81vAjahrib+eNfycl3RRlODH2xd1WWlmM2bUueoS8NTFYIv+qJ9st04oDe2Q/RIvuGV
JNk/hoxUuaLIcyozQvnwX0nrtJzelgu351Nz37TERqXBWNl/17Z0xXize6vkNotwa72+PRr824vE
8rl/XwkvZG8cOCvedyUE29LFz/Fvo+jKKzSkzZr1+aoyAK4dM7FGyWUgA+i5xS8dlvimYLcEXYxj
Nf58r4uI0TOOXkjvihH17UvpEWCNRsMWglnxQtrxkvK8wQq+Q9MtIfoLVrF2PzG85bj1KgTeU9Ez
1JquOI4yYwq7Rq1ADsfgpKGkexhFsRkjm+Bz8fspJWJzc3MDjeUPLiF1BHcXNjsF3jkHJEpMxErH
u59rTsoPgTCLpBiLZzAvnubE+qSjAitDSCT8tFaj9mEongT72TNY850iIbV4oSwv34r2xA0gG4Mw
jy9m5VLbLg+Rmxb/atNyrLJp9dLDQkoY92uMYz+pZJ3ojHMopdv1WtuoMKnA+25aB///uWz1yLFq
smkqEK2nYA3Y13o8wduzxYwmAql2fHZLDXfaF0orKP7sS0p47FPYGxFfESzUwc56n4j8kdquhG6A
CzE5LCl2epEKwuKtGw7AEqKeANv5rfJDPZJwIPa/wMhadRGQWwC8WWccrHNylDTCD7ogLUI2a/TR
EbEDg1G3n75UJs2tDk09X0aIMpCSxr/hICuHo6/X4Tvsb/Im1YQoNB4UdpYxdEovsWkd/mAgw6qc
u9IaPbTGU7S7bSCIPjFYDWoLqj4qa0Jb52iyuoViFqpiaDV6WelOXBcyqotDTyJ/wef6py1KPzas
JGCl8gD51boZGeeOSMfAx63fwAueU7Z1RfueghxX3R8zJ/8EcOSN4LoSCIQwtY1SjBFaMcWRHnyS
QSPI3lC5yB6VUkHxwe4kVJ3G9pzmAFkM7h4qQ1Snh/tg/xTHmQot2fORfpDPMk7kZqqVJEd7PAwN
yI4baLbrjdSOXfXeBli2uP/Vr5R5k9wkRhKwrxCQDCo5C8YlsTHvc5LoQ+Fza5MHn794e2NyRpSs
GA2sDfoj7oXKd5c4XEDn97iDYfy+OhG8IZcDfRj3Ft0KoFpvO+iD0T1BM3T2ob0IMVi5v8++OjoT
RV1951XDilqPjBpAeOB3Kf667oSW9A7ZaiYZ7LFoFSjEKr155C1CkpGAUbDOsYBDV+42U5PH7315
vpetlpFYzI/WJszwE5jG5zQLHJF6gUM9IIF4s2DyniABFkzmNfj+aZbByB85/fJ0ANQ3ZmfbSXcU
5OcMPhWxmkLVIedSskKQRzs6jo4VFPk/KEAMzyZ4CilcUySF4bPa/+nbzjzmFC+2FvlLXXDMlgrT
Anvqfk2yv5m/cjk+iVI2XR1kge/4YztVc8iCgkhCopQCSk8V95hBhiqeTqwf5cVbBHI7OoBzvQep
FAS4U5Fl7YW60uWjAoeRCRCIFSpiOcA92cw/jgxuamvIPYAEGAZ6kce5v0qZ39eABOVXFVpmdd1n
LcODe0eKkGF2UK848JRwjZEsvHUqU2hKkTOzt6Hn7LSD+KbYN4+BTtmmfWZSxIqa/rfpVccrykYG
dwPtP4boR42w75RKkePG0BLqGA4n+k/scp+sClyp5lWMp3PHI0j+yDMwSCewMmbAjglNgzVo18QJ
nYNhzUPkGVWLAWYtagUNjDYbffugVypWRPy9AzopjrBpvRIq9IGHHu8K4qnQwCVMOQjmaffpyNwr
4813mMWL5PKOK/VsoQN5ETrkOzbewdeKKDrcCGQUqcbJd4nqvlTTBYxmVC0mk3lGl0EjllaUHMyz
pEC+WrkJrXd9Vt+bou6lXPUYf+b9V1FyhH2Fkxvxt2iAij51ZS2dmY2Upe6zlS7RhZEnVY+7EIkZ
YxucDO1oJuCODE1a6BzihMSIJjYDZTYZyXeFjlhU08wU3LoBzIH2Pq0CqxqlxVDQyB5qG2hUlU3t
Yr1GmI0zpWBmdZXtADgaWQkPYUm27bwxyAw8fcaYXRj5DIx4EUM1r9qBD+/tza1wqxYoneQoVOem
CVogAeiTPCAzgDQd6r6MHh6B1A14lulyA/1yZfMrhbsxXgMrZ7NHzdhsVCK13aflg55Ag0OAHStl
9cnciMgbJIjilyxTPNKrysm3py1qyRJKXR1N5FwxML8X5aCqsZsLav1PTZBWIvcW4xp7WPqwmCWf
W3QxRoz/MyoileQbVyOi4ORBlNu39+yV/ImixBtEP3cSs/Nhi+gr14WtmQycRiOm+rg6sdBfcZyi
X7SyruqXxm+Hkm0GXcNLRYMraoxEw620kOCBYeTjmcb/3rXnnDyY8csDjlzZ9cE2xDMYMoi4o5/k
I29EUiJlxRkkawCZx8jxsAFQ9s2qBf1ORph5+4OspsH1hXx4o0ytRGjQyOMCrvNiMw/LwJXYt/TU
Yh5+PmONeJhvE+9Txt1eG7JfAqUNIFw6hhNjvreIQSsGtURRI8vxqn9Eb4VYH2/xparpcTwoMdkm
CxwgfZK5WfggLooBQpquy4ghHb05owePGhMZMUO0U+n7WlF4ywCNiDFP8fCy+7EyCPKqTcBSYB5o
efVFyGJ7wCPpsyWSXc4Y5r6dCdCLNCiaiwB1brc6ygz2uAcfyAk1b/Cw70s1Te+Oiz9SLfHYfody
WJq0BgjFaxHWR8tgHuTpuwe9PHzZVFbfxYW2RDgHzN4QUjmDUbR/pXRX27/dAJB2XGy0X1EY+ol8
CGyO8FhJwyYbXJJjeaCCHvFGCMbjXr2O+ZVkX859j1+uLDdMKCvRlBjaVJbH2fH0+SQvYxfVokY4
S/rBsl2IZW03NtahmfgL1K8lKqguloxYsX5gtTYGzr3lb9KXljgzVtkU/ibtzl13cLxOCi/ePBfE
iFgwVBAA+nHgYLH7Yj8YxIC8+FB7G+kPZ33jwg59XiOirccz7kF2tDdvTYIGUvHZ/YUWoVSUnaOq
wG2/w9InR7uGGNjqz/86byUOGVoxOQ33g+txlDKmgDSn2F45uK6ylvjdgIfgxVdy1nM8QkboPkoq
a1x47wreWO5WclzMtXAlDzk5SH4aXpH3U5uWwiv6L3anjuXsa942iZDhwV6saoxqaB9wxbNx6kEx
9Va/CeqR4RmrHwEVBOFnJWfiHzdH0X0YWjMVKRhYwT6w9BcIT+Od+QOZnpqVR6gEe3ws/K1ZfyD7
uHTeB/LVchup+95cj5Ncsl8yZrCCcYaL1jC0o/L8MjWoYpXWBgB6I2r/xoCGJbJ1uSjPpOJc9Vv5
a7Ha4zV9tUTjtztjsK8k65ubAlpYtK/yZeEzalG7kUUufddoDs85aTDR+IieaaeCxhhOULjEYCy0
BvCFXCzSnYx3Gi517amC52HIinZ2jX4GSZb4Jo3u1czkKPj/AYSZi0yt02A8fiNn+M4BjVSBAUkW
uqcIv/lpdZBmba0QyVy3F1a4QUZVYb0fyXZ8AgEjSqUhbS39685ws+ZqxdVNr0i5l1rynWxtKj5K
ywDgNXQMXOzfCfVfSL7QmDtwkY9GP+moZvSC+XdSiYu1zyF3vXOZWMNm1sq0ECWWubBue27pvr7G
nYNiGDseYpmcWS7ewDgb/GBy+fvNJxlnqfrlLKjurphiG2/Rhi9+UF0pk9t5FsB6HpCsNNrk7oTn
9xdPk5M87j8WsA1vvk5KMp0gou18j0++hkVJ0iudcx5pv5MEeagckjNxstWU77nWNSysjEMl/ckg
zyIfxDnqlILyc4PtR95b+PdXmMLlfrBZpp0XuYqtGVa42p46+meTbsgtE3YJrugv/iMN70zlCk9+
q/STVmETJuoCI3u2VBe71uZ0rEnr8rfmWkFh+mMIh5vNi6vbNxNVJpfl2sDUWCQCPCK0x5518QXG
FsOE9e/KtHcR1jdumu/lLDLWiJMCwE2yVPsehdKCPV9p+byM2l3kZI6zbAGmT1Z4x/D29MKsQCfu
x0UXAkrr5c2kZpE4E/+5Ucfbb9dgfWVmTW2X4aKQ5cXTEY7A7pFgpuDPE3B8WzdJMBItN3woQEIg
9T1xVUH9AuAOpxvKJepw8d86WNAhaqtw8ah63julnLSZem134ut61PNBDO+oUhwjHLuE4Sh0OVuN
LKekeyzQC0RAovQn8H6i1RE22d9wNc8B46ztQNmPaKtCTaRq9eNguTY3oYMNxHShalHx4VZ7xByz
vA45vS5f+gHNEjS442Rx+clneWgMw36RKqOHdfCEvjmMhP0xi846KvvcfedxD+JnWr5FK4MlZaAs
iIxfvbDLQyNNCoFjsVneGDn9+tBVntncs916JmpY2/Cukf73q06sz6fRyPnAMmmAe4aXBg9YnVMF
foAtSwdbLRlod53VuGudhmNRXWv6PLjYUKSd+gI6+fvIyMQ0JgPrVXBfXi3TtpYxWrnXn2NXCNoF
djesIXmC8zafnDU6tJDP5CKnPQP4RgYzUK5sLSsIezH0Jmg0GKvVy0UFfUALxIbLL/ynvQ01WYvl
Sz/77mTAKl9OyB45G3gG4AIXm0P8frmifLiKKn4luWFaLoILgXgQX+Y5CZJFQjg30cUDQbnpejZT
s0/EpWmO0BipCK/B09kb6F3Mw8oqhq1MvtPZ1YC/hJ/dWl6G0lwoAAKEDaLTfkT0mV1rufxCb6KR
c1aB6+UEzuT6kY95JcOT3O1Dn12HWwj6rj43eHxk5I8Q2IgQVzZ+Rym7u1Nwuv4NdyTpDFj8wdWl
muwhbcPsOqe5c5IQ7sDYIhygWV8M2cgtOzm/g6I1Zgzu9CBeHiC8ax8G8vxjG4K91f6M4rQTlfXG
O++CH8yi/qD7gPUPPdKfK0Q2CPZmmQ3H1gRpfZtcujXQxwgJUvB/P3ecc4vJsjD2YqZGtDnb0MbP
xVV34bfqaXzUFX3D4D2jlPCIRo1gEZwxwFWvs7yikxojqUS+O3h7Hcp5E8QRu5D8IWelr+AFw+08
XJTh81cyNKWbkExD9nlKBU+nPMgpsWWIUaI9S+RSB44NqPFVmR1ORODfzD0e2VEKNEdcgsnKhpZC
RR+KkqtDIztH7O+y2rPiChL35oFFFy3PR5707HyM+1dYqqYjwJcWQqcBx3PttT0rDqw9uJatc8Q9
QBI/Ia+qm43HJvwkmnd96LzVHgNNorMLooCxwndTuZZkFgNPwmZQxyVie0szvu6fYWuK5WYWtW7l
EFDetsesOwBeWq2CusFn3DKllaDNTHohYLVv+mWY4q/ODoOX4lQmZxjQO+jeO+zMBvYVhi1OMBvi
nmrpagUO/hhbacc8TgfoepoSsZ0l5OJBDvtPns7EQa/5EhzHaWx6AdN2JMTrGUR3fj4J5aVOCqbG
k3Q7kpV9mxI6egOuVfwACJFTkSyMbm+EzhhbYp6FBHQOfEQbHOzh1itCI9QTsvUC6JEOAHRF9xxp
DUI5kn1mQSMxVPtzAfvpbw/JmBwIB4Y75WnP9/4IdiQGgufcUqCSY7DirmFWmpOHAnAA8h+YBvNp
XuHWqsYVH/21zNSSyH5hbzfZy0tXRemK1Q8formuorqbvbWrzcwzSAzS7x7gNohlHHUAeWJ2NZeE
28D6bGcensH2hP9/kBl5gXqz/1MS5imn8g4yZTrqTVleJGAYnAscvmsz1O3P9AuUBM4zPaI+MGlM
VjEm43D+W3Qec57OdHhGcbpqMwzyu/yOoQmnJm1akCz/cbmZYon85l2O3Eq1INJwwoxmehlYo42R
PnhpRbJMLQ74iZ+8kDE5wn7YfYmh8u9UnkmNZxlmzje3Sq2jG37wHgc7KnIXwOvxBiW1dnBe/8Hk
AlKis5bkBX11IdNs276fMXGzfuiY9yPojSpLByQJkqp4CARypsuj6QtI+4ReJiuQOCzWIeyH7mzH
+W79eJGCjZq5SlmfrYa+RMZzONYIDm5jV1Ulle2PFE7avWbC17g6EyL/7WawJbzEGeeKit67u8t6
rr9xwcsQxtbf0PJcgxVxqL9170s/X6TaTwtF94rsDoXkYvBkpq3gC87FEcODD5TEfwJwerbKWiRY
eR4pRys8OrTD1QI4mJO+zz8C70BU0rWCAxcC46tgHjSUXU2YBs2gyC3+Fosdyw+yfjJ8zNM/GFld
iDrPVnO7eIsSLj3q7A+cK4gL1THT5pkhOLXeNBhXHBQr5z/h6z7bTNf4uketR6pYJt+h8NquRtzW
LVlC4l2YgLx3bfk7e2uqIc44Di6do5OKAxgDrEmXk4qwRVtNJPBw1qQ9WaBF9QqXPEUemF9Zqoat
6rl7Pu6Q97cH9dx62kg1c6zKCckj4n+t2JZoK2BSK3xlSGJTeP+raw8wCVhCzknDbEf8bICvOj/2
lKCC2OWpRotGeB81kOue9ziYwM36vnGHUvQX/aJDe9A4jx4Cx07sDY8CniIm5lwi7GzYn89J65A4
gYeW4rocyEXzZUuZRJ6ds+85F46TfavxNwk9SZ6//HS1xsqE3ov/xoN59lYLs2DGjak6c3hcayaj
+j4fiF0RgSKIJGnfaC8dTKhdynYH/6mtmXI7PgRgVee8NLUzcn30JMD4lTPkfPN9+kKBIhw/rPGx
iwZWyfdsfX1OyIzs9YPISWla2FEhJXqGZ0OT9MC4pijN83g/Ex6SSeeClOZKszLjKzTsg8Nj6NDn
Pt3dcrflPgN92rUMXa1ph4XiXFm5vOUg5ZjPY4hyGK/4Wb5hPbFEm09CsJLKUHK/z35jx4Ra3yuw
J1o0e+QELcP2D+LKS5LtAHJOqXvc/I7TiQRv7jCUSbGZZnArKlv+WWESXskLvWG0yT7mtdFLbGzF
RTCqPwCB/nBKXFZJ4pudekAXoiZArxc5V93S0eritiP8+oqmLFt/g1+pR0cmeYH5WUvrPUJXZrSF
Lcmfr3ODgvB1uCpkOMivNkeWqa7xnMQ4/1C4VgWQo97UG9MtJ4hntGTGSPHFJAJKSrUD1/4wWDP5
28nRgu0l5tR4tSynMM5SwhJs93KRenb1+Wh8Gl+nOYIoSOP5WfX2SVddX8culcpCU7uyjMauxdb8
aFKhEWV/DBL8vDmQFxdORCBR762ytxT0DzprMzcNKMu0XYQ1K0Qj+NUe4Ij9/g4oLVsHEcXvjSbS
mNjPpm2rNay8z7aC6Dp1yjjVNnEF8Jl626MQyqWFfSCJRm1gdzyNbUqtU48RLWNCOrLdF9/b8ek2
c3f8+ngis8jCh+2I/RlLy+iWi7lmzv+o/qE/YJUX8TnXemju05A0RmOnr/DGwI6xCJRDvyiRI24v
31DeRM/q/twQRQzuA0piMrHj4XAtqLtqHpqu1wRdcYE16kkD40mhLwjEBJYCVp/HOR6icqZhwOPJ
lfgmgeSCt/Mnf3t9aE3Niv71rx1CH5DstUwUwS2kuDLxmEg/IYEd6vnktSEK+RHThhiWS1FeSVzv
nBEEKI6p0w7tggeLzzOU3aY9K324nXRE8fq9H9QyiWuZQB51Di/g2SmgjdkXLqTO1idloDmbuO8Q
4zWptxmkWI4o2SRUH61kL3wpZDf/WbeR3t+szXHF7jR7GJtLA124G44zXYUBWs/I3ib0X0ww9cg+
a+AnVRi9ktbDSqtPhDcY+pxYNlaFChQY+LuVOu/+LAoeCk3WGUkWu5AF4Q6B4rSCcUHgQ7KtsrJ+
4UQ+4nWUsd5n77LbWXXlrSK2NxpVacN5xoWqG8cGIx72IDdxan1m3yQVcLFBfEa4y2Ffi4w/kl34
bndVX2ids5STvRqbGf9jkq9Q7hY4n4sVTi9Tco3wcQDj32HFNYabnYd+0/qIUD+D6Jvten1i1uQP
p8TfrfkV3/rBvaLGSqcqwfpyh1p1Jb9fm4eIh/DSHBLkbwBOo2JRV0E+VkNXnnZwIjzIZYNEHg6A
Ss8tFiuebfj4bEVHg+iap0AcBWzOv8aUYILOKVoLBFpjdl6kThNgioX2oVVrpX7F/4w/QpVSQqRG
w0ZpPq90DLDjp+ryRAqIf0PrtlP+KmpZpGQ8JYo29AqIxX/jn24I6hxQxRUvyDEwzNx2LkM2xM7u
K1J9/wBoXX1l3s1JeLf8M1aKQAzZofBuiFgQeW+HEnGF/gAO+tACaFDGpJYBTYsa1k1yF8jxmPyk
nDpYxCr7KkRrnwXLMeRn4m8ryB3rcOI9J6rzJs0zijfPWptRkheLiM+qxygXtw00M3PN6dv5J2C9
TenkCCqpoMCNReda/oNxP9GBGrmet1jfL5fKspfsHWI0AWL2lpVUjstLOU01JerJoRpRjdTptgmW
jUibK2X6OT57/H+n3TcM4tAp5pF4RcExAJ1qjmFCAHloI4YoU4fEuhQ77jerXh27K0fWBpN0tWRZ
QQYpomh9rasYDKP0LNwNkq1E0SfnmI7Ib+wFcM8Apo8UjKhhrCEaHZ6EVX5e+MhK8nwMjLAe4I3R
X9hkhXXZzV9Ang9fFync6igTFQq1PplVoxjQMihNcuywfv0KnWLRIiv4QtxBaIO8oJNS0cbAcLlj
L6Q+n2tOimOfOyGxDJsRwHgcj0pVAEPlejb5iOwHjDWmTxHjMDoY5J3XacgSQ2pZA3GkAsiYNq8G
LReAna3k0C9aNQFx7u0s4WjGFtLFhHGwCGNQNBf1SHEDpqVBTW7W5h2QvTbs1bvqGwAsILktuL71
DQEFfrk602Bxu8BsbkJq4hfnDufuk1r1BN6WaB9IQreKN5biFCaJang3k1Kc9DRnWiv1NWwlrA0b
SQrSCYvi2VrD9auliaMwwgTlwOiuJF7DWrTzK6xD8o00SsL7XatE41QeTemZHIz48ftN/uKCX5JC
q8V6M7k2EZCbMHF1OtisM6lVHmAHNydgeFCmZ2gfVhW5/56RyIfSvaHvjRz4LmuT+j/SSkfrTvty
SKZ1s/qiJ1GJ1dQywD5LLGHq6sPDFI5jRD0aiQz/5i+qRRa60gMgfdtyRCP0YoyyX5FLwp1ZBaIg
OdmYaCEV/HdeljW51rXrUVAJmGKwZN4phg/CULCT9e0rEM/eFnWUKB42BPIFgy0CPbWP7hpo8tn4
eB+LKeCuMRXi+gb417L99/yZOuxXsp8baVxCSRgFwisjaIKgrAItXIX/pedU4bRERt2GnwOW72H1
oRcSbCnnj1apbikUan7BG1L8Ciuy05A4ObFG07H7tF2Op0rR8WXK6Kz9OLdXuzFEcJdD/mxTgMaO
ybtv4lkbcjQxJGaR2QgNoeIxS4IKDQUjMVzjbfsu5wK/lZ/P9E8TxvDP5M3kmXWXNsdvFOQloR9r
quxbMw8zdmXLtKC5hRQaHmCM/LFDhpneRquTchWtGzjkt/2/tknUmBf/NaZa7eH6xlYk2oj8DZ0W
rC62ioRMSNEnhEJm4v2PXDBBqbvaM1lnpPfCCz0BV2q61mLgyCEvKAxsm+/vPNwOZsh/tE0eF0s5
FF6h4DMG72fjmBFHlyHd0lY31DQ9TgJ/MDP20lEYME2s4O8Xi1V5nVSU84zbJai8Ow+0tYVRbb+m
B7/tzFBArxf6MU5b4vWxaSdITqCPcGyVEJYtA1pWVMDNukSCQOqz7Y9liT3PAY1E6Kj65fQs7M2u
2qHdID6YS3YbyzyDD6dwenC12Sl45/AIWIwNOGCW161j7e/z63sjMtH3gghXQEH3M3UJxp9w+F4G
ON5AZ/MKl1kZ0wtSo/7TVjnsG3nK5Kb0GYbBwX+lDFITliqOI3Rv1KOgxgIjd3Ouh5CaCINSfpFV
1wF5ktXV46ct1J4Xse42QVzCEJFaDJdjBNOQaEcot2rzndkGafIAYX2f85MtsU3JZV9mVmwcEBsR
WHlg/7/9FJ/Li7F44pgWU8/SmfL0OWRgSHX5SbPXh+VHniPP9YDIzoMkHt+AxklKof+4uqm2Lf9d
tFTBN4cAbPIKg5opVRl5mSLxWvLdWlVG5GraQCfjeL1SHLIRl2xLnRVjmFqdlsRyhm29Vf4ZjrIC
CaiXhWia4iaWZ9vKd7nQQD/gyKAd2v8nGwm3+SqcMM6bZV+EQ1Oiq1Lg3T1k2IzJxWRnGXFviKro
xeb7mkGaPUg3fSIMpMfBw5NiICw/APH/nfH/x+qxi0NJnCsRmr6iXcoGCJ0erX6t1fMmUBI8pwjJ
OwJRyh93F9JlwP0nrkEmT47AeCoT++NRY02McJ2ACJGS99sCCxgf5mFON3SLYdUdiIKWvnPXna6J
qx8+q1TxufXZurppvbJgVXJB0IUcNyWQT2b8KzXHoIEjIAsgX/HRgKKVz7z1uwG7cqKhNfgdVmLg
BCEzGPTzfj/F9bPXDh07IS/eFdtT/HmWZvaXmLlHKiu6kIzD7kwkxLv5kqrABwSU9scw8z1FXLFX
NkfFzGsVDFztuXOaHYC4dmIp/4RrfrozG6lT66XUZvXNncwDf3HjvqnviuEzA0HM7ti5mxSOrRtQ
JrEsikTCSaTlxGIZu0xTgV4fFX1rjwaKJhnR3Uj8LTmwFW/tRhGf7fXHHsW8gj8aZc9QPg3O4U+R
l3dQj6iP+O+0boHoqoIGz6zkhGDE3e6SOl2XXQVYQzGZZ8/YKgWKHT9zBLt9YOqG39q+7wXaFWfb
HshGOnH7F9WYvrTDNFw+xjdEqcHWLJ9SqrMGZtLsjDU0+dK6a6v87q2zmO5NgwS4P2gik9UsHk6z
q04n9G97siOi3br0+y1m95hgW1TKvpVepxwLjHDHcQav9jH1jEO6NmkWzcjZ4yBVahRjcPDMt4DC
abl+Eaey0EenrycT5IAUoziqvdPGaiypXRNSVOKku6i0moFQozFDrUKI8dD6fr7VswwdD2X1DtdR
6Q7qCYzF7MaM+zHsq1K2zMNZ7xZ/H9SwnkgfCV6F7e4tMLKIIn+w78ef6b5Huy4JDQBlT2PwPDXE
KDXXzbfZVZVpz9skJFDgQ+5m2AqOchOPHDkQkI76FDD6XBldrDAGCV//iwu2ta9lLRALpC6v4zPA
mxLs0RSOnpNWCRnKOXc7dcdZx0S/FyJueqd+VsfVoSA8wR5IvW4/JQ149bUwta/yXolq7ZvG9CAT
RhU2Oa8soULLiyo39khZU8PK+f6EzC0E1DO51VOKfPBuq9gfLSvw0NT+WnR2r+pypfYCpPbcLI6R
VA7IjUbkRIyUe/R1HIk9CIibNoXvlmzYfr0gBwbO2imflE4HB7lZ/t7zgitvzxNZmpJAcBQBxQsv
U2qVl9e+Yy1saxAbx8DLLXUgEWHaW9xZhucgoCOSLCNXM6fcJjmLa7pMVmhk8wZVsjt8L/FRniIQ
TnUOsvJsoA/z1zEMAj8TucNZbdDsxd6d1byvZGAP19UVPZSlGBH1S+/hiL0xH3qgBkP26FZvoCBM
lzEJbXvAj2oRyZtIpqmAUbLVAOn7Du3oQk6WomW26hXkotKQyMBjYowDZbSjfXAaoiefOy1FTYdk
iTPQBDeOf8haiN4Oo2s2UxRVKxVbIfHF0wj1R1UYZ/HIqTDIJp2STTxCMrHFQGGf4PJj07A/6ivk
qHMjPwe0hKR0j8xlEEPGfqiwyMYkR00WbBHRracb4Iv2v2AJ3NldS0IS7VK4AaAz+8mkZFmrPbGk
euobDd6vNMuAB5OOXh4f558nnGDm5LMuM45kquB2dNwYNw8lkh7zZuVlHPvJMuDW7rRDBsP9dRFU
abLAaVPD4T2f9JUPa4qye9Fcm3XCjDFkOL2RbFakxMP2uBklcuExMK0J7kpyN773eGhN8ilw/AmL
WW2eyf5XS8a8IK77KVICy0smyP6ArMP1dAgDzHGwBfvWk0NuIHpZzR5GwAeduL+cJMg/2xytjXZ5
JQHw5KUR3xiVgVwy+IOycBZJ9tSEGYOxBAfqpgeov+tknj7o7kFfdRhdYdV7xWSjZYESvc5rZtUA
I1UU6bPQCmymzmP7AVFzPp+I6faT/+psJXc25x3SlWxzhv62G4L3ErBGDlxWwNKZgoTZPdtAoY3G
/KWfYTPeoYCbVbHuRUCwTe0oO0zVWSX9+q0Pxe5nvluY9m97FzKgSnTG9CoAlvhD9yQ5g3Tao9DB
JqrW7MlrPb36Y/lr6BCHoK+qmsrOW6+Pn4PX4+His2IKrYtIu5eopcG1Z1g8oFqC3fzRWn3eowtB
HTTWsyn+Jw43isfrk8uoT6frbjxrs4etKFoG2erRH3yC9T/qjqsv+YRxgPvXKxlnuyXoY/1jd5WR
7cDg/n2SPhFnaSSYXo2DrKv0OKa23s1xygXfKogJE9AP4Y7DSkFknpv5FqNdh0TpgxAIqG3u6DuU
rSaT3QpSdckhUvm0Ln17m4210AcKBxfAUr6vcZ6mtwBz0MUYIu0XnEUJ/BVp4IPXKyBvR1QiOqEB
Ezx1xZzSjLxBLBc/h5+qnIhIdjjFWEYb6ZnYZ0y3TKuvLh7PBvG4TPkqcl19MXh0sYpeTLuHhcE9
yIpiS2dcv0VUQNfXKJHV6gnNgNL/n1+XYtxfiv/t0ivDq1D/lTCC4RvgX4mIeeYw1dla/sewbMCc
7YGYXeURiRhFwpDAlkVVgMHotiffQNkySkY5/EA/BdMRAXtkLeoZ4od7t5pzURL5P05pEr0AcXxL
5P35ZlCU5NU+gEv1D5LgXhOdpDp9HsvSZst+2OPfJcFfr7a+4lk/yCB3K3N2Or0Pu6oR4qBxT/iU
98yAYKCnAEykNLU+ggrp6PKbmb2KIiES1ar6ds4Pn4DqNIJnTpf3ixyir7buARUyp/RRUHSXkwGy
v4OESBfZ/NsHBMXnJCNLUfJAxZIy6EznyWSf4ly0eK7xJWDeY3R4Z/3GqCFnuWZa/bpnGzmFu7sp
iZaDABiaJhaZ1bz52mgobhP4gJIIOznTPXF475kP4G10iLAEs6pn0IV0AQvQnm0+W3Pt0lhd3QbC
CGaL0xcf5JUj3H6+0usqamA+jzySn2zS4kS594TGbhdw9DPvdWcHbTfi+GqHdlsOl1r95m8amKw2
cLDydPBMD9c5/Hb0F4IEWKDfH25ww259M2zJn7zruWgCcd/lDYb14Ok2vBuoWENrYPmFtmbUMx5G
+IwD3VCSLRUzP7W8B3fYAu9Tssi5nImBeDoT4zDyRA3LmzL7DZR9h+JeKo+2ILnU/V8qjT3DT8dX
bpAHe7JqR2WmqByP4V2tGTKcTmtJdONu+YLPbp9UhvDwawU60Ktrjahij9a3czHXSekOWI5bs9yt
5kYB6VgBZOosOT++AjtCrDhizr690sJHBvT0LNBORqqHrsrVc3iPZvicCiUvArxeKL1dZIxRhEuS
C1y46rlot6cH/2wRXuCQsINkVT3Eb9bFQ49oW25095Cu5rWLhMyTxDLTKNq63tRd4OIEgaPQBuld
NEard/oy2/jrCXcuOhb/9uCqYmneQTHiqn5Q9WdQIoZXJ2gUwDZH8z1aJoC8b8mrpMEhbBl9Rw1o
Alm78JgXQrag/98pOVRZ72T56mtL9xKZ39B97FuFLbZ1b+hZmghGurVryTBweqHPLtDhyzclQ9hR
7Ab3kmPxPiNpMrWiiLOxuGE5GNh3uILvuNUvNJ+Drb4Dt+ou9n19WykGdM7ZKYbexZEJlhpTM5Cs
owypla+3NQqUi2q/C9YtcltQGvPkoZMlmqTne1h359cNoGAz+sKlAjdtW4UnnTgU2scFtTTqQbQI
hQNu18DytP7tbzB99RjNyxd58botumbJn3WtnFv8jdwOd+2BgObVDNGXLPh/5AFLsdcbi9c2uFtZ
79ekW47YZrB8qaMIGllZC2ZQotVy3+Rpx6aS8GJBflsgNLE9DKVCWt3W/lFtIJWmoY7Ak9yZPQWq
q0qxMMRZ5mvsTyV5gdNV+T+GmFZGAg1VnnsTgRR5WmebzHcncEAaKqEWG1wIQOOVcwMGzwVN7li1
bPZ7tFBjgNVF0abE1bF8Ngam33gCxei6SIof/pEzzULxQiCrAFzQhrOykRzhWc2W99PhDZnqudzv
5HXwUuyoTfHQsUBwW/Z1urqOGv3+mcIb65Kd4LsG37DeJM846PyGRtUv1oC4/eIxeLdvycomZ6Eu
SawafT94qdTfql04QFGk7QLrQ1VNjuC5RbV7ffNQ20Cq17t4Em3QPQrZqRMXWNG9veiQT9QZBRxJ
TLrFRmFjqfLrIOpwv0Ta/+gXA0AejX7TFZMSwcL/qV4BLOhSBRckYIGYpwwaZdVpMW39JGS1/RoQ
/2hNwfKufii0k+NQyFtQXzI/zypnqaiHpGQF3LOq9pR01/ac5lYv5Kmhxz/B7G6/OA8mFMret4bQ
fxEyMU7O9v0luYB17IgPOlYFiOv3HXqljMSSDcy+OWpFK4P5mqCgk2vHVk9hGCEHGa1r0iHGUha3
6K6XXExg46gYccXc3tlkaRap9aPzSEbvIcL4KcU54QUSgG4BqDBJh8aLkONPzqfY9/QnOpLH3MLC
U1zBkEJ0k48KXeQocVZSRIW4yFY1S1IR/A3nMNnHRdYW6WB6J/kxnw11/bPd+jJ1Z1U0ju1cbVkD
SkDM9+Y+tkjkPfDJQYoEqlzp9C5bDCsqW/QHevD3+OewGdBf7y0r1fznrlyBpje5UF27s7QKlzwm
5WRYCYjjprUQGA/BuLUvbhElr96FqLiDwPToLD7fLuDY0pnIeTNG6kDrozOhmKuykWIPJYIAzrpo
jf7b6m82WOGfUOysUenCALU08Yqddv+FNAjGeOkKF+wCMBVpI0Ah23q3yah0NgLLyXDbwwSaAoVu
+E+p4zqfg1FoKQB5RFx2bOOLHtDWZ+WMC4VOdG1YIUZkB0xNEGxzyIC9Edf3DNxTElUSfkUvSPSL
q3V9WkaTPqBTJP7qY5YjBYUoGqzdEMC1GPduhzQyZRr3UAuDaQEtMQsmjkEM2yFqoho2yja3/Zyu
WydkLeg+IQnz8BwtYwXNRiLfJUGf5YzuEanEjuZ0h86F01Fe5v7zou4I7El/cu7YI7XmL/MoNZrU
mJJTEeP33MjRUduy5zjZsOz5dbf16hEiMdlmycbfoFGnp0wnk53rVBA38a9hvobRHK32ktrd9ulp
BN72Bo2Rj7xBX0sAiBs0MxgvW8WcCCcY3gpW4jLFb5XhAR0E88JS25h0ICkIM6nCXQcSWNuG2PIv
Ys0P5+1lidhW3mREKFJ6KVtB38cjKFIn9Awv19jRF1oS9d0Bi6TY5T5hBFMmnFLJv0UsbQ6yEWSc
Oe/jgbG2rONDd0O7+5vMSFikhFxL3+PFcvIaMcU/InitRvQ1hpRe/KBxGa9bhijTMmT31tCBbGdj
FYEfOmSkvJr94i9GT6nRvBatGDBlUumXnH6x4M1qsMtfd+pmttZFyG2gZYGSpfpUCBbcj7fBCy7M
+LAfBqgM/Miog2KcyyyHI2M7P9HUdc1Zcv7Z/paFVawGLojQGlIi/Mp4EhdtVRdYrYlNNf04Fy8p
E3HIVHl8moCMnF7LsRAVYlQ11LdCD5RMWWT7hw1RvUjruu/nsgBPPNSqWsvwOlvelCwvKyIKSWrl
HJ4JBtS3zlrF5ITDeKdk1YVJEDEXGMF6z1C92KEwfVkgc0LAwHNrztmK6aB7lkMfoL2A3/de6ATK
H1tyF3IpeuSmaFHSnOfUq5mo8zQEwOKkEyCDoO6HbE3Ucr8nmS7KFZ0T48NksPbgoWSpGAMKWm0A
SwO2+6QA4dDI/B46flGTI0fJ9wrii+XUJtFlYeAnnV7aq5KyMRIF5PhU4CgJ5MQpmx+1RWaEom9f
au6a+ZiY+SlXa/YZbix78oUmPVbMnu1qpre+/q81qujDZFsZjvaAm3ocyoPct8epTeXAjSLF6kWL
FeVP7GMP0BhTWR/Z0t5Zx3qssG7pocs7WAw5mdYBnZBH5kEGXuD5GX3EBulzU2zEMfP+WkY5ygrk
EA/vrLU9TzLX15EY4OS7xllaxMDJmzJZD5Vv+HNSqYvbnb9eRLt7MGTX0bhSazMiTkZUeLr+QuiX
ZHH47fvPUh1fd94J1iMIWDXAcVucoaclA7dpXCd1Y3OUWxIFpG44Itettk6PZNK5s6Z7E/liqRba
jeeq+VzzOptmTzsCaA7JcY3dR6o7yEXKFQG9Zdi67AfUDThvdarU+x2GMZ/abhPLbdse09fRPm/N
mvRT2AuuGF0GXPAz3l7YaD/jWG5GE1XHoBF3sbHWeZiownnp6UCPyrdcaJtaUxYP8IoNqfEzkn82
PMfLR/Z2mpfFxSqgpCcWYwUZXfIYU9vxL6HevMxWc+zfludov9lJ8SgxkMVEKrmd2CqkYpUOsUzu
HVFRaTLfZj551cH02Xfuj+jLzpvi5yQODgwfr9+NIaiGWGmxORW1MqjhsFdgr7u/40+femDTWZZn
G8NqLOafsaWjd1BNjs5mk9kOjJKC50Kd+ZznKkH1RPIQX6vUKbIPtwtZEAqJF6i1dtLhtirKLu6K
D4Iy1BKQ2RlC/rPy83UsZ66umI6jbs3yhlP36wb2TlSbUeV0FshdTQ9QzKJqvzcx49/bGyAWAHpu
JUfQDhGsRQeNSo6nuTKHIumF5aEO6j2+QKAVzGRCyXLRK6rLTvuG9qOh4fuQmjCnGzoQNsvo+pAq
tRa3x2wj2JHflyve2DZjVwG0YSSP3XXpfcbl6JkR6cNQY5xDDIHdMbQg4DXr/aYB/Rh2FkBRrtNh
fSnys1SWy3u5IuGL1QUdtPY/WOm7e5OaWaoVmIBSuHLj2knDUc6P3OfnmtkYBXX+R4nkYm74/7Wq
R8WYteg0VtIAxMznQ8NHkYDW+1+bNf1qYnOAbiAMwpZTUCmdL8j/tEzb9y/vKPAX44QrWkhW/oGA
MoxiOcPO/t8ICYUDjIbN+ytvPr4mL0+YqDmXBoxc6bILFHydjTqS4Q2jV3xj95Mh34ySmqQucqJP
Zl+rRknX1w9+XrCpispfR1dUIxAVRHxy234HuFZF0P1js8u40+Fdw1FVh7G6tTJ2jMgs36ng6s4B
juMwgk0/W6+J8ykm4yWMoGRBcyjR828o/qHTpEb8NclpPQH4vV6p6PZyXtX5ljJKJs5fCykG3SOz
wQAG0YkuBslhDh1WlSP/q9dXSj7w5U5OB/8zBU7GEh20+E/HA5Yg2pRZUFiW1Du0PwgG0B5elvXC
LehinoZDZGC4ZwBS+npsGuo+cEQ0/lIY3al1Ao426MT0QBRZGjumuwiczUJ6MvUWQ3eRlTZ40l8s
dIP1b0Lu2fqxDhmrSTtf5+oUEDaSs8ReokoET8606VGBWpEp1FusAEaYmuBjDFGWRWUNBuNkuskN
SSrAoWtpeaQwa7qwUIcYY1dqtBCKJ5A7WDlEu8vRni0VreZJxod8BpwDEmsfgCnPnUivODFLT9xY
mxIXPP8mIf9zUlzJ2Ca5hHmGLZ97Ng+Y7oCv/nAzGpcLf61kAZKDxx2H5W5ysQQ1oAUEr6kWmOUR
zXUJ6RKwySndkuehLBS10Xoc+/ZUQj2nBXJR9ZNQZiarSaV52uOCAumklc3MIj/7eLNLq3o/AH9C
a1uAkPdKLD1ADtQRyz7UwhAk5mT//2hxBoS/YzPTtTcxE4QN8PK4cLtu7n2Gmk3wZ4UVVnYJPhhj
aEZHNkrT6Xll0zXMbIKIAn5LxsUJ6KKZ7dig5J4V5F9yMVQojbnRPvlbI0cD1BNOYRwoUt/Wj9/P
ks4KPBsqwi3Z30r6m6Kgo6gHpooB8zyXAsfOwPR94b2Eopyw6Xi1KT6cbOUF8GGvZtMJhjzsbk9t
eFxVCyCC8U4Y7uddi4MX0zyTPTL6bjWi1+tbkgpjbPV3Mrhff9jX5HimBwURuETBQZkwpdlUcDo2
pMT4BZjQQEOeCwsPBZHtcpAJevAuhJKg0AlR9wpbUYatoMCflTRqe4WFmqk1sFt0xFpHktTatE8U
JccqQ7hV1Z+jTPQ9c8m5AQHwkT8easAtlMk+rDaaXbYlrX92rRjFKsqh/t6dmLH7HeYzDeLjmaxP
vx353sGrZZ33EicSKeK+/BxffK6J5gCbDqj1BKgqH1bi8T2m3bsNTmMgaF8mQOXorBKoW207FCdK
7d2YGv+Vr2XILJJUgzdGaVjKNknezCChsR/FOuRTWHBB0qHjXXd9T6g2QfkBMeGKrOm3K+Wb6Gwr
th5d6BQ5Img7UmWd1qmGbYoqaJj3z8dxMEOXBVxaYt8Em53pfaG8XT3Ax4nwKxunrJgQsZ97/X43
2LMFAGc+Ut2f8QoKv05hIGpkId5Xm0kH5+wZRFOWgw1UNBrzeuAngbgaPjD38gRKjzep7AXXb3d6
CYoftb9ywI72BOWeYgAj/kvH7JKInZpICs6AhMFrjfD2M7GOK1J1sl7Dt8MMAdIDCXWDz19WLxrq
n1P+Q3GJAC+GZIYCwR5qiZLbWXE+LrhuOkPwvXnSiNE35oF+rYynqvNxmzKFQmWUgPtzWeR62Slc
xb5Z+9+ZMvqyPJLGczJLqx/RyQAFUG/qa3Yec0NA3K4Wdtmvnd5LeQbSNN3pUMqXLICyQzHNEpgD
y7jjcadN8kEn1Hv1P7RwlPR+66FBeWhdBXQ8fv/O+cazdO3S14wbLl721mswQwY+geOqQgsVeVPV
snfO+ptNdz7YdknYCUC57sGTbiY4eCGq18r06xN8XXQ1BV4Y0FPzhsZFd8moS7KnSPSeD8plDuEE
zdYQ10Ax4lQ5JEHnbeOKU49xTYmVN8P8OWKjJ/yG14+1wwrUvjD7Ff5ICksJFP2QXgsYCxGPl7hg
Q/rbLxjPG9A6yl8NWzl4AkbfgZ3+gBuV62UlUKQjkAdv2JRQmSUoZrUugpS0GgNE4QUHmhfhBMGX
6REnG5zG9jh0wnmVzPUXl+okPUPDul/btXNyrPen7SrVjUWkdRcc9F3x6p+IInJIw5jaG6HYrEC2
a6dVS4MxyZndgM70rvUwtClwMCzDBusP9plLSkypEzJF9yhpb0l93A6v0boTtOFMPzHxFLSmPFCW
jI72uvBa3DBa2GoWtK0HcGnXdfk8KLokS5sfYIu8CIle/II9jWc0S48AGrICqEpd0M4Mv/o15xu+
kfrWebKYjm0v8XYUdrtHr1ohOm1w9dG8iRoJKjoLKlXYzIwqR1Nb8lpi4h/DQBsXm6p+21TFTWEH
ij2M3in5XA5qgESuXTm/KS9vdLVTRVsR4eSa/k3ARLJHhqMV//gzUkGraiqkxKTRoTA11NYRp6r4
N+k6wxWAw4ZwVyCoKhCxAfO8W3zF8835M0+527/IraxtJN1rtDJLnrZ0+tFTfz+5VNawj4cs8XsX
6NmbA2ox9YZLmy+2pNzCDYi/vGQihRC5k2JNdwWYODubmgYYkF2JvTuHD+vOQDVUYAxh0W4DkGMy
JVq+dGL5OgXJbDVbipGEsTK5bNJf1PK5y7irrfVdoyt6/TDR0+wHk+uMh1L2G44gIhzfJVqQXvl6
Ai/1wM3kWHSOdz/ZFlBUjlesg6Am05TowC95Ya+Ynv7OAUFSO/OHmXvKKUdCZEVkRqFpnCg411V9
3MHQ05oJsNuYdLaRV0n3H8poi34FCrezDBK+DnFhwRv3HAuucyds21zvTREaqR1BCTlbV8v1h+GW
p66U3/Mr5Pg2SSJYaeWH0uiSJTsCxLlwnZYhni9OYT2w2gUCYq1MmY777dIQjnpA3udYmk3+fDCP
xlC2pX3FHdhSTzMQAYAEr+lgezF84poAlTfSiPnQ8bkx7WEDYmN9Ar9FN5ZYmYE8ufUHU2VdT495
4COy3nL/GHQm64le1WdQd1qirm0awL784NC7OMmkZNJKFG6GyJlHPHYc4II8cDBgpUWKFwgJ1272
D/H8aR9kPuyexwe95IqareKCFtP739DNGRB8jw0r9dl2Xa21L+F3dJhKsAbp3/pjq2zgbAGkzZya
GqWfOEdzAuVOELkbGyo+1Y6gVQbIVI56M+k3zQol/scNh+vMbisFhNHf2Dfkqrnnd1UnFIFK68F+
rEMTND0MTnK/f/+5yQnMIepq0N23E4/zePhAPAj1ZKu7GzsYJ8YXXdw1foyJyTSoBXtFPTHadKYC
/SmpdVGEWI3f8BS/wobpJupEvMoxQtQW2wdmHOK8p+a7fF56cpu0IJHTzqS/q0urgldlekQw7fnV
cxehWsBAKvZkoL+2PTtfxx9vfjxvflFekxlnhEYfPYm9WTY7YWyUhhQUqJu2r2rJ6HjMj6IkN6jJ
t3RoP388Rmo985/GIQmrnZ7R9Yuyqz9NA885pFAyc+bV8oH66+ScqivvBMVOMZ36cZmejHDK0UJ6
nnxuGED/8zGhmN6fMgLy0eu2jcwbvKS9FNtk39baWDLuYKQnCOETzgkBURlbMaTp+sQtmbUSJzV4
QysqyuH7baJJvKTbJxQ0HmdulW5VAGy66buD7fNMNEh6nzQOUprYZlKw8te4wVIpVTO6s9VprL1x
HhtJOl1AVaYsTgy7SZTlIbhLswQ0gPuK7zDfWEFiDR5Zeh0xLNPY9yBjonvXPGwzgrCLI0Ltgmt1
gn+qqRyZQjSCOn/7sr9G0MhetWQcTx8MtRV9+bDZRoHkW6mO6/IzLgk8IjzhYO1koYPNsrIdCNcj
SrHjEkYFz319uGym9vwszEBi2DnCnLo+iCLdpqcsOobBn+L0l6UTUIgbXYDxmwO1HnzXM1M+dfDx
TGVSnRjg5CgOW/afaDUA1d6W/75RT+HtVlFbVk1fN0RxqzdrIg0tsw6kr3VOs/v+bYAEQoRo3wS5
ZnrI5qrFvbkYQ8cGsIZPt0Z643h4iethrdakd6blXTvJ1tO6Zu0EDxfRLqdAr4ai54zG1tsLAcBY
II4/cuWNkXYT92S+Ewx7MCsFner95IjPASQK3pQZaweYvLqpDcnQOMEHSp1td7uVyLxjq3LVf5n9
kLbJRVLiZYT3/cOT6x3IDfb6lPVafnyQ11uiy+jGmU7n44DEdMHqjcNVfTsgByyozHlxoRjcAaZ+
D+Oj03ehIyXEhtR9stBY83Elv/b/Sv6CE0gE/TfvTxwyiAJ6M5+Jbm6f1+SycHiKjvBr0cmtAMEL
JsCQpMLMn+k1AavNwm5rQ0iDsFNRj3902NTff8dMknP4B860SyoLw9jYQeqvpOananPLPV+3kV02
AX8zG0l/15CZGDjTsNoSFaJma7WKTwZFABBTzn2OAPOA6YqqSTvMGGB/5FE6wVhHGFU1wO6QDBsM
pF6D2A+eKLInE2q6NpXC+Ie17mUZbsuhgZyWilPxULebH+DERK57Sue7RBM8ZCsryROIWmQl+Di8
rpY1nPGXG2GPdpGT85MoxVvvzupxJFVX9++syY39hvZHCljuj/XlIraG7g23ccIGP6sHEpDPXFqX
SWXgiO56ZkpA856vGhCEkJnmXLalwWjKXVDTcKDEQBW73vFDtm7DwdX1Ry9p/+6xDbuCSyU9FTUs
n1iGInlF/uXofg9DnWhCCSKTSJrBxYi7m5STh5qRbKPRVbQCrsBR5aBS0wMDMkLQa22ziKf3qwOF
un5buGtJ/Nf0pDK4B5/+zVcGbD335OSAhtliFFXocBzyvnTxpcfmMcokqcYlibiNA3TJtnEZzewj
euj8xTt96eqHI1uX7KZw7XcRPSq0GCJpy80YalfUMOP9OgQUUKtpmO3+SgcTLOKV9/1tJKJIsC73
ZViOPvhqo6eVfgGBSL8Xb28+HIJf1wNdp2sBI7W6Y05kz3vHvZx4tzb6ZkFoQCm+rgFOTuz+FrA4
TUmiNDea5GvB+ZYRF4zrGZXF6Be7B8rApjNCaXuDpD/uzcVCjrITXnOTT8KvjHn8ikuVUBzRBg69
umgzanUdntnQGpC4Ea57KYi7nbjTPoW/mnSKegqs/vnSysN6K9hb6+f/ZlP13ECzU5aPqcjSumSV
9Mfh9ZFmD0Y4IuiNLh+VmBch7kWO9KMM0fX4D0GPMe2c4haYdF8Dkd0utjDfdI38AEvwIPJTYZJS
bmQbvk9HnGCL3HBTUMHYZ0dVb9b0JjyoG1/eolRqTmPyIb8oVVSUHTDfUSGO4Ia32A9dcx7Fn8J3
8FwJeghCPGVY4bEDcgHxlIZTJe+EZMJh9Ds0QK69zktOp7QOZkyOcO2iYvcCee3vqBAxvfU5GE6b
nPdLKVlSRxcS7kvJbPUo+hxx/M30XQ9wK2xF1JQLgKdHf2ewtnz+c7ioBpzGpryN0V0VxD7mRfam
NFs0zPcu6B90UL0gjXduFMMMABOQw5hCCaedbTtXsUishirqNG8R9T6jqw8OAW/00dEw06JBAQ37
7qCoNkI1EUMvKVTD+vClAzuZG5+Nic1+HJ8W5IBiJdzEja3WQZNJzqX16W/spFIBgWLsz1GrqM/e
4W2uVk3dO4ZmFe7Z1R3h/z1x2vZvHD9dYeNWDaRw600/q86PsWyryZLdle+eI1G2dHf4Z1uyzJ+k
yzc5qOICpZHTLPRnYttngo4YmSytNLFEvBpQI5vo3gckHSbwMow2Djdf6nqmvxo019K3hUtAibfy
v8xp+Dof4kWQkzwXZQTWVn4Pahz9LsNwtC7nHx++TYhT3RCxxBxWTwM8kojB4Tb4BfddWby6OujF
pKe9cwPZAWJZfBjUPcfX23UDSypBCagkoA4C3YJwrUXh5arsE5RhcQR5CdhcWeukG8Jkv56ftRpP
bd+hYkE5j3S8Ggxys+iG6zVbrIEtRCcxU2dVIqB16paFgywKO1IK0d0ohcvwUFxlqYVPlUvrINhE
ukJbRnik1906d95yVHRMgiUOU5rT/nCEsrV/VQgU26otaqhw0mF5FBu5Ns3u90cMuJ8YS7P0QuUd
xScWSu9FkAExUBZVsb0xm8QRKGKDOv3nr4uf0JllNe3TACD6PtJnDGt8SSETa4fIIxPzy3I/9XMO
1J2u+08q7jOL2KDGErzx65rRjro42GlgajfHmcMJX8jxjJlFioHd2PG372H+Pij+X9FCDO49zKHg
jWkLHwUrJuQIe7KJrKDl82GA8TpoZOnvnDL+H01f9zEcJhU/Lop4IOGdwtC8XNUlQAqgN/R2rPiI
9QaxXzuSiq9+oLOHxuuYbxgKtUC1PpR9YKd+nQvna2+LYu7w54Oux01xEeOhPnGu1ntVWWcrZXk1
2PSAsGNNVhpZyVhky0mzDGCnpnzvDsFXKVaVeC7BiIbdiJucSkVc7z6OllrjLTkk7QGz8V5CK4Qq
bOa0JVXmj2NODNuyC14dsxF/s7JKXBmmdTwHoKjcn5UIT8MEc1rFYqSo+g9p/2w70E05T/MAIYCo
Igck0HGf3T1qz1lcVOI1MxieAEBAGX3Khsrf1ev165PvaaUyJNPOhL+ktWYxGE5/hs2DElw+h9pC
LWGjJouMhx/FLNxB203oVHiZZCSGHt2HrWh2Rctiqv6nWPx7HJ8peOA/NGdOIsE7F7N3FyHItOI0
fPwdRvCwMZMSviVkKy76F8GbGnhxWyHmzpni8k9ZtMVQfjEgAOmf5wddnYPr7QngCgz0aBcfy+IU
NnD/H4RiiHN8DSZmyHV6IieYYWNTLMqEv1eJP+y09ITeRfzoMIDAWshiPvSrhfJaUo7/0+Ce6jV4
SL8NOlo8cIRO1mB0ogS9zFAAf+dEizWqUYWrhtPa9eIccBT5KEDa8seIOgVm5d/fAZb4X6u+2+4F
biMOgM+MdASj0KZNbl9ktJksCYABjU4QN4yr/DbHDGZWrgzgMxtE462DmKN3yY6K1NdOH0QmRiMl
rbJKYjJfUMuoLAb3laSEeYYm/vfW4bFPOZ/OLiQXcddD2KTg3fb2lthxhVRTvHYliWLUBXdxrr0M
X+2/JfqtdwHhRcz4+bOwBjc2LrnDinAkreDZciNuJ6HQR36R8kAYXmDWWMxIAPOokYotHhb3sNIb
W7wXGndl63yrOsnZUGZX19UfFGH6z8ftg8Pb9mfRUst2vUDcohBK8HV5fZkpJU69FTjs8W8BIehL
nfaaktyjd8DRz213f3iVkSoEZHjVTINk1/Utrq8jXoC/KfuyO6AfwKSL++pBPGwlDyw7TrTaufDe
M19DUxqRebpeyJue4ntSM/1nj06AdOx7YUNkQ5ejhbOk5o1fMG5vA5gncKpzxEdK1Q1CQhsK94mg
Ojff/ADtmB2rM7swnd0acdNV68RyrxjMykR/was7xdKd0Tl51lGocUS/GKzSWOVqKjy355TNCEES
X7jZGm74INuQhMYD1Y6qxPH5TmMuljTxySgowyBOtLQhC7+Ii01UJSpszPReNZDipWZRpBR1uvxz
hjsZzuKzPJbSktTtUgMrjwgL4HP391bZIHRrZhe6s2EUVvEjyh6bdQyM3DcfczWgRiuh9HinPYLl
l/M8icrisMNqIeWHfCtrdDprJXpypww1cpErSWZRKYYhd8yVN5MX7OalnnxTrS54epgsIvUtOKjf
LBLFM4d7ph+YPYiotbb4/zqQ5dk7rRXIia7Hlp5iZW141kGD4p8sUBgbbCw+K4X/At8qe6K4PnV0
a/+LAjzq/1ylwIg9Twk9XAlzsIqfvAHgagCdqszgWtHZTCQ0bIb1Z5I+fBNXJvksT1miN30Irce8
6Vb5BxDE9VTAOb3QawfiMK1dIPpM5Ww+l5izTNZDyJxQqNz1i3eUEi1+oP88+sRiHeiR8Tq7GInY
5pSvH5IGuFYib7mX38ZYB5W/Y6C+Dz9G+n8MvoJji2g0bMv3q5nlW00JnGTPoPZU1BpaRqu6yAM2
llAIZoCW3yq58s9CNWhc6SVKUAIEHVtI8YL7hf8lws0fzp+bRkzAMGNk6KbiYnPaPoRprirZg/KL
w747XHwQPvR8YfKt05V6wt7DZc9VvXAe7AL60BySWH3hgZQdISBz6dZebHc40RiOroTbpZSWOCmH
ybVjD0UO4UPoMgJbCHYVDQge2iLfC671XVKCtXUUlL2Xwxp7BUPR36yly/J3RbBVbftTpmuPU3Qa
HC4XcNXuFv6y02cOKd3Vx2dXvVYVI5dfwrhSO1Yrvw2VQBLcLaWVcrh8QZlYMQn+ZiKZ3wQ1duQp
Vq2Pze5tqehsCZVCKlcJEXgF/F9dDMiHrnINJaMeEcx50Lkk+76vOr2VB71BxigkHrLSEfvl+ab4
ha900WvcU51aFdfHQg27+vl2U/oTYZubaNnqpNAgwtfHbKiY5/boszmXDrMtQM7w+z5o6OtjeJR6
mrxlJgfoe3iWlOMEVPtnAMohFhNkesJP3by4YWjm+8TOgt+t6zHI9nU7wh8D0dJ3vd3rb+2EDkFI
AJy0WUsJovkoR8kmuCz3F0NFOX3rGKcQB5Q23pi2PeFKW9Yz7atLiAG1jpYkazMKv8w9Cn29sddY
R+TrIJdOGUl4fBFJyH6nwOsVVhL4Mf8uT7uASp7Jc1UwWUn+Oojeh8YjN3egdUillpesZe48NaXh
IG2B0/gM4E8jvZhowJdGrsk+IOpMTZLPrzslfqvJbB2h35pCa8CcCnaxo+6ymSxpCK3eyED7UPjl
MPD/40Qk59QcQAyGF4hcVTIfS8Sf6s5qe6mejG13R9EzkDzvXPH59bqe+bzncw5jHCJwcmqhFRMI
xbMz5i26yCVPnnNrMJpLA0F7EOphiGt+gfiYQXFJg5PCyhDOCYi6ARfqsdjI0sWRYabdyYSK6pwx
AGvOd8Sd5zhApuQdDyxiBbhTDLnMh+8+9VVtQlv3h5wnoh/3KGcxfLbPdJgmGpuaTbGnuwsnkR6b
MVb9XcMXxlhjERHYef71TU2//t8f4nDJgl0SCHmSe8qgcAYcJrOk7Y7VdJZ5zJAn737YycknD8L7
yxAt1IULuTHBJEORg575Fq1zr7XGLQ5dlbyn39SrhOmBuhdPvhUMNCZNwfQkjKXrTt3hki4mh6uK
K9gbg2t8DDncHhqnMjPQ4agh8/F5smXxIGbNgXXn3Vbj7Rz/Qry1Nd9CKqZ6R+jFoss/rexydmtJ
ntWKopRhBjmjqLyFGCa0uiPgXaHsuyFydSQGMm/GqQdkBJej0B8xe/RMfDbu73M49BY0DAU+K4rL
/llFGGu0zeKA/RV2mHIt+5iS+gDfQA2VAR5LWICGoSFH+9EVcw1fXhNH8p5jK0A89pn2V3+vCrUb
r4ZMCME4BkRWqKUmlc//Y/sKskmq3bCscZh1b7NdEXi3yBgpKKU1bW+etS0F0FT/YuK5H7CcHqyi
61A3FAapZNESG8isYa7sGcmGjh+I3NGUuwszFSRqlAW2ZfYGhBPInPz9nRQ9AdV8KM8Le67yYFeC
+jmjJFMQAOUXskTwCcGH7mkyNO8CJdL3bOressvFH6VIdYbshPhLrD2fVy+oA1GUILa98T3Ig9de
GZvUSbkjS8fb928jMTn9I1pwNnwzQcYDnzD/nJ2oIdBxV3P2Bv2h4I+/g/B3Qy2hNdi2uywedth6
w2qBCAlFrclICug2tTnd9wzqWlDxeZ2qRTTkBGC0m0cH27EUvXKZvP8NoT3bYuRl0WEOy4NcTZdR
zak78XEOiUwhUMwUG2PlGM2Se5AzUr0esIh6mrVb3Uyzyf84oA5W/GVDAU98WRNEuk4Edx/B9F1L
eqbUz+yQeZJamQKku/Y/VmoZe8uBWQWbfcgG1Vxz4RJ9UpIaZ+SiUC6+A3OXCCti/4A99GyF3vNy
CDEXi9ALLNXM65S7Y99oc1QgCQOaetQ0ovM9rc7IvRAhSmRlfpn5HifxWqac5QRZXzcNlys5O+F/
tvfl4CYB1RtF/w8I1HCgLDd96dhYN+heZopFiB/7bmmssHHIBjxiTNViVyQVLW09b7S0uXt9y+N0
UnRTsfIA0oJOB6l0JVb3l4d5D2ZKRviy0mWsOkOu5URxSXFUj/aYaNvAwJ+ZlwGVkKS51XI82iJW
VgBXkxC1oDnmrgbbzsOycqTdwxQeOhutmYyYRdwryG3saAcWzfmJ/ex9vNLPc/NTlFTa5r3z6Glj
alDjGY+Ii8753py88r7+nd+6U4ldoitvCCHK9zUHN9NtPt4eoiYVn/8f/5Greyog/uxQ9p/VzL89
AKWmdjwUvyKoHw/gs9OoFQ25JBPbiffEL4wW2x/S/WsGfxevETObo22zoYE7uw1jAu23mbDgkzZp
amMykwgFYcIvl8sApa2yjUw3N316oI///KWHC2mbOJg0HndE2Jiz1wVgHk52tqg1HgBRfp4tf1Xg
Jp2LoeIR62bHS/SXS2GLGVS3cT0K3KdOvYcfK9NtbqanNsEX7FoC4BXHtAAiMlH9L5aFCKLcAQSF
TyBcHVxHzeffaDDFAqf0VZryQb4sTlaCRFKOub0BVzdY30S3iuESkpHlTy4X9CltZtJ+bVJ3VcCb
2/W3mOktbwPe9RYPucN7KLiEJS1LWiYy2kUEkgD12Nmlv7fEx24o3DuFjeBEiisXDdiJQtgwrA7O
co9j+W8Z9COxZQgwSon/UQTFaC0vYWida3K+TXTZdgde3i74gg1ewqQ1+UToeNN3TjUgwWwNJ/3O
LYrc50TDM4OZbTp+O5cHCpQZM5LBtk4Pha/y8fYmLphzeDvPIJ7pEz3FDj5B7amEpGXe1ewbia9/
GRtu0V0dJ/lv9tooXwvVpRVS6VLbL4UBny61W5gzP1f5oN0xx3HtVZH6mCnheMrmYb+cXct805rq
7NtZY+WERT3cjssHMRE62mXQm87gXWHXg2nzloNsBNkWniXeyJutG8H8QsFgHlRfS9iSuIEZwXlq
6ZawiOdx1NGCDjT+DhPNEXKc8aJKubx7ZuEDSEehJQ/Nl2dx2cGtrVxyWleCk5UThAVJPoc70H1b
1Z5iybUp+mLhIlPknsYVzvwBqcd/ol23PGI6Z8NoHLX0ANHBkPU/1ARsdKxkn/4A+lEptMNl3R3G
D63YjgcTYSHGpw0gKhmCN2viLqnHFXOA+tSFTIs23bliuTebGd2wTZ2DM2OCk2QLL+/0HJs5dsRE
2xKw1bQJeqTul6tJE2EUU5j1PxTMrkq3ftYYOhJu9t9BR/+/XpaJR+mnfjiNzGZ7EKkcPNgKGwz1
9NJ7hin5sP50vWwcgbVCWWmSxl4Kdr1OsjpeCSIc1vkLoZU54LWaBBJh9f4ywQkrkDx7/q7kmvOH
HMWUo/fLp2fRZxw/ttZsQJUz8UrEuR6yB7yAA+DepIMY43SNDaJ98qXwNVNtgYAJmyJqmT4aEMOb
/3Fc1sfySG+iGFXMDr5dp2ui/MnQkwYu0nGLzTN4maBZ0Fc82VhY4FzPtTQlP4hVsQ6+P2XPjbjq
lW8A3RSHrBnzEL7Jx2a3Pz+j/nJLAbWBO3NN6P7r3B3r3+TnoOUQNlRD/fQIfCA80fCzn8GEf9m8
qlJQUvzjrOAkcutRG1vDzQqS8Bs+khwlbiUJ5jg/K4/y6KQnwUP2ku+96S9WJpZ3wGsfjvfzW2Ob
eIWkh++kTlCWKon5mV3Sym33wzOEsXEjAa0QJHrn0b+MuYtUCOwVpCF5Ol93OcGicxjFVj6Kz6Sx
dIQ28cQstQSigKUELD6EXXMmFYCM4D/3isINbQuEv62Rkx77Tn+MZhP6BfFDbNB/DodoUmuqIgyQ
Eup3sejG9JlU
`protect end_protected

